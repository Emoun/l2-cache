module Rx(
  input        clock,
  input        reset,
  input        io_rxd,
  input        io_channel_ready,
  output       io_channel_valid,
  output [7:0] io_channel_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  rxReg_REG; // @[Uart.scala 76:30]
  reg  rxReg; // @[Uart.scala 76:22]
  reg [7:0] shiftReg; // @[Uart.scala 78:25]
  reg [19:0] cntReg; // @[Uart.scala 79:23]
  reg [3:0] bitsReg; // @[Uart.scala 80:24]
  reg  valReg; // @[Uart.scala 81:23]
  wire [19:0] _cntReg_T_1 = cntReg - 20'h1; // @[Uart.scala 84:22]
  wire [7:0] _shiftReg_T_1 = {rxReg,shiftReg[7:1]}; // @[Cat.scala 33:92]
  wire [3:0] _bitsReg_T_1 = bitsReg - 4'h1; // @[Uart.scala 88:24]
  wire  _GEN_0 = bitsReg == 4'h1 | valReg; // @[Uart.scala 90:27 91:14 81:23]
  assign io_channel_valid = valReg; // @[Uart.scala 103:20]
  assign io_channel_bits = shiftReg; // @[Uart.scala 102:19]
  always @(posedge clock) begin
    rxReg_REG <= reset | io_rxd; // @[Uart.scala 76:{30,30,30}]
    rxReg <= reset | rxReg_REG; // @[Uart.scala 76:{22,22,22}]
    if (reset) begin // @[Uart.scala 78:25]
      shiftReg <= 8'h0; // @[Uart.scala 78:25]
    end else if (!(cntReg != 20'h0)) begin // @[Uart.scala 83:24]
      if (bitsReg != 4'h0) begin // @[Uart.scala 85:31]
        shiftReg <= _shiftReg_T_1; // @[Uart.scala 87:14]
      end
    end
    if (reset) begin // @[Uart.scala 79:23]
      cntReg <= 20'h0; // @[Uart.scala 79:23]
    end else if (cntReg != 20'h0) begin // @[Uart.scala 83:24]
      cntReg <= _cntReg_T_1; // @[Uart.scala 84:12]
    end else if (bitsReg != 4'h0) begin // @[Uart.scala 85:31]
      cntReg <= 20'h1b1; // @[Uart.scala 86:12]
    end else if (~rxReg) begin // @[Uart.scala 93:29]
      cntReg <= 20'h28a; // @[Uart.scala 94:12]
    end
    if (reset) begin // @[Uart.scala 80:24]
      bitsReg <= 4'h0; // @[Uart.scala 80:24]
    end else if (!(cntReg != 20'h0)) begin // @[Uart.scala 83:24]
      if (bitsReg != 4'h0) begin // @[Uart.scala 85:31]
        bitsReg <= _bitsReg_T_1; // @[Uart.scala 88:13]
      end else if (~rxReg) begin // @[Uart.scala 93:29]
        bitsReg <= 4'h8; // @[Uart.scala 95:13]
      end
    end
    if (reset) begin // @[Uart.scala 81:23]
      valReg <= 1'h0; // @[Uart.scala 81:23]
    end else if (valReg & io_channel_ready) begin // @[Uart.scala 98:36]
      valReg <= 1'h0; // @[Uart.scala 99:12]
    end else if (!(cntReg != 20'h0)) begin // @[Uart.scala 83:24]
      if (bitsReg != 4'h0) begin // @[Uart.scala 85:31]
        valReg <= _GEN_0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rxReg_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rxReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shiftReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  cntReg = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  bitsReg = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  valReg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Buffer(
  input        clock,
  input        reset,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  stateReg; // @[Uart.scala 116:25]
  reg [7:0] dataReg; // @[Uart.scala 117:24]
  wire  _io_in_ready_T = ~stateReg; // @[Uart.scala 119:27]
  wire  _GEN_1 = io_in_valid | stateReg; // @[Uart.scala 123:23 125:16 116:25]
  assign io_in_ready = ~stateReg; // @[Uart.scala 119:27]
  assign io_out_valid = stateReg; // @[Uart.scala 120:28]
  assign io_out_bits = dataReg; // @[Uart.scala 132:15]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 116:25]
      stateReg <= 1'h0; // @[Uart.scala 116:25]
    end else if (_io_in_ready_T) begin // @[Uart.scala 122:28]
      stateReg <= _GEN_1;
    end else if (io_out_ready) begin // @[Uart.scala 128:24]
      stateReg <= 1'h0; // @[Uart.scala 129:16]
    end
    if (reset) begin // @[Uart.scala 117:24]
      dataReg <= 8'h0; // @[Uart.scala 117:24]
    end else if (_io_in_ready_T) begin // @[Uart.scala 122:28]
      if (io_in_valid) begin // @[Uart.scala 123:23]
        dataReg <= io_in_bits; // @[Uart.scala 124:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BufferedRx(
  input        clock,
  input        reset,
  input        io_rxd,
  input        io_channel_ready,
  output       io_channel_valid,
  output [7:0] io_channel_bits
);
  wire  rx_clock; // @[CacheRequestController.scala 13:18]
  wire  rx_reset; // @[CacheRequestController.scala 13:18]
  wire  rx_io_rxd; // @[CacheRequestController.scala 13:18]
  wire  rx_io_channel_ready; // @[CacheRequestController.scala 13:18]
  wire  rx_io_channel_valid; // @[CacheRequestController.scala 13:18]
  wire [7:0] rx_io_channel_bits; // @[CacheRequestController.scala 13:18]
  wire  buf__clock; // @[CacheRequestController.scala 14:19]
  wire  buf__reset; // @[CacheRequestController.scala 14:19]
  wire  buf__io_in_ready; // @[CacheRequestController.scala 14:19]
  wire  buf__io_in_valid; // @[CacheRequestController.scala 14:19]
  wire [7:0] buf__io_in_bits; // @[CacheRequestController.scala 14:19]
  wire  buf__io_out_ready; // @[CacheRequestController.scala 14:19]
  wire  buf__io_out_valid; // @[CacheRequestController.scala 14:19]
  wire [7:0] buf__io_out_bits; // @[CacheRequestController.scala 14:19]
  Rx rx ( // @[CacheRequestController.scala 13:18]
    .clock(rx_clock),
    .reset(rx_reset),
    .io_rxd(rx_io_rxd),
    .io_channel_ready(rx_io_channel_ready),
    .io_channel_valid(rx_io_channel_valid),
    .io_channel_bits(rx_io_channel_bits)
  );
  Buffer buf_ ( // @[CacheRequestController.scala 14:19]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_in_ready(buf__io_in_ready),
    .io_in_valid(buf__io_in_valid),
    .io_in_bits(buf__io_in_bits),
    .io_out_ready(buf__io_out_ready),
    .io_out_valid(buf__io_out_valid),
    .io_out_bits(buf__io_out_bits)
  );
  assign io_channel_valid = buf__io_out_valid; // @[CacheRequestController.scala 17:14]
  assign io_channel_bits = buf__io_out_bits; // @[CacheRequestController.scala 17:14]
  assign rx_clock = clock;
  assign rx_reset = reset;
  assign rx_io_rxd = io_rxd; // @[CacheRequestController.scala 18:13]
  assign rx_io_channel_ready = buf__io_in_ready; // @[CacheRequestController.scala 16:13]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_in_valid = rx_io_channel_valid; // @[CacheRequestController.scala 16:13]
  assign buf__io_in_bits = rx_io_channel_bits; // @[CacheRequestController.scala 16:13]
  assign buf__io_out_ready = io_channel_ready; // @[CacheRequestController.scala 17:14]
endmodule
module Tx(
  input        clock,
  input        reset,
  output       io_txd,
  output       io_channel_ready,
  input        io_channel_valid,
  input  [7:0] io_channel_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [10:0] shiftReg; // @[Uart.scala 30:25]
  reg [19:0] cntReg; // @[Uart.scala 31:23]
  reg [3:0] bitsReg; // @[Uart.scala 32:24]
  wire  _io_channel_ready_T = cntReg == 20'h0; // @[Uart.scala 34:31]
  wire [9:0] shift = shiftReg[10:1]; // @[Uart.scala 41:28]
  wire [10:0] _shiftReg_T_1 = {1'h1,shift}; // @[Cat.scala 33:92]
  wire [3:0] _bitsReg_T_1 = bitsReg - 4'h1; // @[Uart.scala 43:26]
  wire [10:0] _shiftReg_T_3 = {2'h3,io_channel_bits,1'h0}; // @[Cat.scala 33:92]
  wire [19:0] _cntReg_T_1 = cntReg - 20'h1; // @[Uart.scala 54:22]
  assign io_txd = shiftReg[0]; // @[Uart.scala 35:21]
  assign io_channel_ready = cntReg == 20'h0 & bitsReg == 4'h0; // @[Uart.scala 34:40]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 30:25]
      shiftReg <= 11'h7ff; // @[Uart.scala 30:25]
    end else if (_io_channel_ready_T) begin // @[Uart.scala 37:24]
      if (bitsReg != 4'h0) begin // @[Uart.scala 40:27]
        shiftReg <= _shiftReg_T_1; // @[Uart.scala 42:16]
      end else if (io_channel_valid) begin // @[Uart.scala 45:30]
        shiftReg <= _shiftReg_T_3; // @[Uart.scala 46:18]
      end else begin
        shiftReg <= 11'h7ff; // @[Uart.scala 49:18]
      end
    end
    if (reset) begin // @[Uart.scala 31:23]
      cntReg <= 20'h0; // @[Uart.scala 31:23]
    end else if (_io_channel_ready_T) begin // @[Uart.scala 37:24]
      cntReg <= 20'h1b1; // @[Uart.scala 39:12]
    end else begin
      cntReg <= _cntReg_T_1; // @[Uart.scala 54:12]
    end
    if (reset) begin // @[Uart.scala 32:24]
      bitsReg <= 4'h0; // @[Uart.scala 32:24]
    end else if (_io_channel_ready_T) begin // @[Uart.scala 37:24]
      if (bitsReg != 4'h0) begin // @[Uart.scala 40:27]
        bitsReg <= _bitsReg_T_1; // @[Uart.scala 43:15]
      end else if (io_channel_valid) begin // @[Uart.scala 45:30]
        bitsReg <= 4'hb; // @[Uart.scala 47:17]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftReg = _RAND_0[10:0];
  _RAND_1 = {1{`RANDOM}};
  cntReg = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  bitsReg = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BufferedTx(
  input        clock,
  input        reset,
  output       io_txd,
  output       io_channel_ready,
  input        io_channel_valid,
  input  [7:0] io_channel_bits
);
  wire  tx_clock; // @[Uart.scala 143:18]
  wire  tx_reset; // @[Uart.scala 143:18]
  wire  tx_io_txd; // @[Uart.scala 143:18]
  wire  tx_io_channel_ready; // @[Uart.scala 143:18]
  wire  tx_io_channel_valid; // @[Uart.scala 143:18]
  wire [7:0] tx_io_channel_bits; // @[Uart.scala 143:18]
  wire  buf__clock; // @[Uart.scala 144:19]
  wire  buf__reset; // @[Uart.scala 144:19]
  wire  buf__io_in_ready; // @[Uart.scala 144:19]
  wire  buf__io_in_valid; // @[Uart.scala 144:19]
  wire [7:0] buf__io_in_bits; // @[Uart.scala 144:19]
  wire  buf__io_out_ready; // @[Uart.scala 144:19]
  wire  buf__io_out_valid; // @[Uart.scala 144:19]
  wire [7:0] buf__io_out_bits; // @[Uart.scala 144:19]
  Tx tx ( // @[Uart.scala 143:18]
    .clock(tx_clock),
    .reset(tx_reset),
    .io_txd(tx_io_txd),
    .io_channel_ready(tx_io_channel_ready),
    .io_channel_valid(tx_io_channel_valid),
    .io_channel_bits(tx_io_channel_bits)
  );
  Buffer buf_ ( // @[Uart.scala 144:19]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_in_ready(buf__io_in_ready),
    .io_in_valid(buf__io_in_valid),
    .io_in_bits(buf__io_in_bits),
    .io_out_ready(buf__io_out_ready),
    .io_out_valid(buf__io_out_valid),
    .io_out_bits(buf__io_out_bits)
  );
  assign io_txd = tx_io_txd; // @[Uart.scala 148:10]
  assign io_channel_ready = buf__io_in_ready; // @[Uart.scala 146:13]
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_channel_valid = buf__io_out_valid; // @[Uart.scala 147:17]
  assign tx_io_channel_bits = buf__io_out_bits; // @[Uart.scala 147:17]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_in_valid = io_channel_valid; // @[Uart.scala 146:13]
  assign buf__io_in_bits = io_channel_bits; // @[Uart.scala 146:13]
  assign buf__io_out_ready = tx_io_channel_ready; // @[Uart.scala 147:17]
endmodule
module Uart(
  input        clock,
  input        reset,
  input        io__rxd,
  output       io__txd,
  input        io__rxChannel_ready,
  output       io__rxChannel_valid,
  output [7:0] io__rxChannel_bits,
  output       io__txChannel_ready,
  input        io__txChannel_valid,
  input  [7:0] io__txChannel_bits
);
  wire  rx_clock; // @[CacheRequestController.scala 29:18]
  wire  rx_reset; // @[CacheRequestController.scala 29:18]
  wire  rx_io_rxd; // @[CacheRequestController.scala 29:18]
  wire  rx_io_channel_ready; // @[CacheRequestController.scala 29:18]
  wire  rx_io_channel_valid; // @[CacheRequestController.scala 29:18]
  wire [7:0] rx_io_channel_bits; // @[CacheRequestController.scala 29:18]
  wire  tx_clock; // @[CacheRequestController.scala 30:18]
  wire  tx_reset; // @[CacheRequestController.scala 30:18]
  wire  tx_io_txd; // @[CacheRequestController.scala 30:18]
  wire  tx_io_channel_ready; // @[CacheRequestController.scala 30:18]
  wire  tx_io_channel_valid; // @[CacheRequestController.scala 30:18]
  wire [7:0] tx_io_channel_bits; // @[CacheRequestController.scala 30:18]
  BufferedRx rx ( // @[CacheRequestController.scala 29:18]
    .clock(rx_clock),
    .reset(rx_reset),
    .io_rxd(rx_io_rxd),
    .io_channel_ready(rx_io_channel_ready),
    .io_channel_valid(rx_io_channel_valid),
    .io_channel_bits(rx_io_channel_bits)
  );
  BufferedTx tx ( // @[CacheRequestController.scala 30:18]
    .clock(tx_clock),
    .reset(tx_reset),
    .io_txd(tx_io_txd),
    .io_channel_ready(tx_io_channel_ready),
    .io_channel_valid(tx_io_channel_valid),
    .io_channel_bits(tx_io_channel_bits)
  );
  assign io__txd = tx_io_txd; // @[CacheRequestController.scala 35:10]
  assign io__rxChannel_valid = rx_io_channel_valid; // @[CacheRequestController.scala 32:16]
  assign io__rxChannel_bits = rx_io_channel_bits; // @[CacheRequestController.scala 32:16]
  assign io__txChannel_ready = tx_io_channel_ready; // @[CacheRequestController.scala 34:17]
  assign rx_clock = clock;
  assign rx_reset = reset;
  assign rx_io_rxd = io__rxd; // @[CacheRequestController.scala 33:13]
  assign rx_io_channel_ready = io__rxChannel_ready; // @[CacheRequestController.scala 32:16]
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_channel_valid = io__txChannel_valid; // @[CacheRequestController.scala 34:17]
  assign tx_io_channel_bits = io__txChannel_bits; // @[CacheRequestController.scala 34:17]
endmodule
module CacheRequestController(
  input          clock,
  input          reset,
  input          io_rxd,
  output         io_txd,
  input          io_cache_coreReqs_0_reqId_ready,
  output         io_cache_coreReqs_0_reqId_valid,
  output [1:0]   io_cache_coreReqs_0_reqId_bits,
  output [14:0]  io_cache_coreReqs_0_addr,
  output         io_cache_coreReqs_0_rw,
  output [127:0] io_cache_coreReqs_0_wData,
  input          io_cache_coreReqs_1_reqId_ready,
  output         io_cache_coreReqs_1_reqId_valid,
  output [1:0]   io_cache_coreReqs_1_reqId_bits,
  output [14:0]  io_cache_coreReqs_1_addr,
  output         io_cache_coreReqs_1_rw,
  output [127:0] io_cache_coreReqs_1_wData,
  input          io_cache_coreReqs_2_reqId_ready,
  output         io_cache_coreReqs_2_reqId_valid,
  output [1:0]   io_cache_coreReqs_2_reqId_bits,
  output [14:0]  io_cache_coreReqs_2_addr,
  output         io_cache_coreReqs_2_rw,
  output [127:0] io_cache_coreReqs_2_wData,
  input          io_cache_coreReqs_3_reqId_ready,
  output         io_cache_coreReqs_3_reqId_valid,
  output [1:0]   io_cache_coreReqs_3_reqId_bits,
  output [14:0]  io_cache_coreReqs_3_addr,
  output         io_cache_coreReqs_3_rw,
  output [127:0] io_cache_coreReqs_3_wData,
  input          io_cache_coreResps_0_reqId_valid,
  input  [1:0]   io_cache_coreResps_0_reqId_bits,
  input  [127:0] io_cache_coreResps_0_rData,
  input          io_cache_coreResps_0_responseStatus,
  input          io_cache_coreResps_1_reqId_valid,
  input  [1:0]   io_cache_coreResps_1_reqId_bits,
  input  [127:0] io_cache_coreResps_1_rData,
  input          io_cache_coreResps_1_responseStatus,
  input          io_cache_coreResps_2_reqId_valid,
  input  [1:0]   io_cache_coreResps_2_reqId_bits,
  input  [127:0] io_cache_coreResps_2_rData,
  input          io_cache_coreResps_2_responseStatus,
  input          io_cache_coreResps_3_reqId_valid,
  input  [1:0]   io_cache_coreResps_3_reqId_bits,
  input  [127:0] io_cache_coreResps_3_rData,
  input          io_cache_coreResps_3_responseStatus
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_REG_INIT
  wire  uart_clock; // @[CacheRequestController.scala 57:20]
  wire  uart_reset; // @[CacheRequestController.scala 57:20]
  wire  uart_io__rxd; // @[CacheRequestController.scala 57:20]
  wire  uart_io__txd; // @[CacheRequestController.scala 57:20]
  wire  uart_io__rxChannel_ready; // @[CacheRequestController.scala 57:20]
  wire  uart_io__rxChannel_valid; // @[CacheRequestController.scala 57:20]
  wire [7:0] uart_io__rxChannel_bits; // @[CacheRequestController.scala 57:20]
  wire  uart_io__txChannel_ready; // @[CacheRequestController.scala 57:20]
  wire  uart_io__txChannel_valid; // @[CacheRequestController.scala 57:20]
  wire [7:0] uart_io__txChannel_bits; // @[CacheRequestController.scala 57:20]
  reg [1:0] stateReg; // @[CacheRequestController.scala 60:25]
  reg [7:0] cmdReg_0; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_1; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_2; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_3; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_4; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_5; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_6; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_7; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_8; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_9; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_10; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_11; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_12; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_13; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_14; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_15; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_16; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_17; // @[CacheRequestController.scala 61:23]
  reg [7:0] cmdReg_18; // @[CacheRequestController.scala 61:23]
  reg [7:0] sendDataReg_0; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_1; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_2; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_3; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_4; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_5; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_6; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_7; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_8; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_9; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_10; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_11; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_12; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_13; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_14; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_15; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_16; // @[CacheRequestController.scala 62:28]
  reg [7:0] sendDataReg_17; // @[CacheRequestController.scala 62:28]
  reg [4:0] cmdRcvCntReg; // @[CacheRequestController.scala 63:29]
  reg [4:0] sendDataCntReg; // @[CacheRequestController.scala 64:31]
  wire [79:0] cmdAsUint_hi = {cmdReg_18,cmdReg_17,cmdReg_16,cmdReg_15,cmdReg_14,cmdReg_13,cmdReg_12,cmdReg_11,cmdReg_10,
    cmdReg_9}; // @[CacheRequestController.scala 73:26]
  wire [151:0] cmdAsUint = {cmdAsUint_hi,cmdReg_8,cmdReg_7,cmdReg_6,cmdReg_5,cmdReg_4,cmdReg_3,cmdReg_2,cmdReg_1,
    cmdReg_0}; // @[CacheRequestController.scala 73:26]
  wire [1:0] rw = cmdAsUint[148:147]; // @[CacheRequestController.scala 74:21]
  wire [1:0] coreId = cmdAsUint[144:143]; // @[CacheRequestController.scala 76:25]
  wire  rxReady = 2'h0 == stateReg; // @[CacheRequestController.scala 80:20]
  wire [4:0] _cmdRcvCntReg_T_1 = cmdRcvCntReg + 5'h1; // @[CacheRequestController.scala 84:38]
  wire [7:0] _cmdReg_cmdRcvCntReg = uart_io__rxChannel_bits; // @[CacheRequestController.scala 85:{30,30}]
  wire  _GEN_42 = 2'h1 == coreId ? io_cache_coreReqs_1_reqId_ready : io_cache_coreReqs_0_reqId_ready; // @[CacheRequestController.scala 95:{51,51}]
  wire  _GEN_43 = 2'h2 == coreId ? io_cache_coreReqs_2_reqId_ready : _GEN_42; // @[CacheRequestController.scala 95:{51,51}]
  wire  _GEN_44 = 2'h3 == coreId ? io_cache_coreReqs_3_reqId_ready : _GEN_43; // @[CacheRequestController.scala 95:{51,51}]
  wire  _GEN_47 = 2'h1 == coreId ? io_cache_coreResps_1_reqId_valid : io_cache_coreResps_0_reqId_valid; // @[CacheRequestController.scala 101:{52,52}]
  wire  _GEN_48 = 2'h2 == coreId ? io_cache_coreResps_2_reqId_valid : _GEN_47; // @[CacheRequestController.scala 101:{52,52}]
  wire  _GEN_49 = 2'h3 == coreId ? io_cache_coreResps_3_reqId_valid : _GEN_48; // @[CacheRequestController.scala 101:{52,52}]
  wire [127:0] _GEN_51 = 2'h1 == coreId ? io_cache_coreResps_1_rData : io_cache_coreResps_0_rData; // @[CacheRequestController.scala 103:{71,71}]
  wire [127:0] _GEN_52 = 2'h2 == coreId ? io_cache_coreResps_2_rData : _GEN_51; // @[CacheRequestController.scala 103:{71,71}]
  wire [127:0] _GEN_53 = 2'h3 == coreId ? io_cache_coreResps_3_rData : _GEN_52; // @[CacheRequestController.scala 103:{71,71}]
  wire  _GEN_55 = 2'h1 == coreId ? io_cache_coreResps_1_responseStatus : io_cache_coreResps_0_responseStatus; // @[Cat.scala 33:{92,92}]
  wire  _GEN_56 = 2'h2 == coreId ? io_cache_coreResps_2_responseStatus : _GEN_55; // @[Cat.scala 33:{92,92}]
  wire  _GEN_57 = 2'h3 == coreId ? io_cache_coreResps_3_responseStatus : _GEN_56; // @[Cat.scala 33:{92,92}]
  wire [1:0] _GEN_59 = 2'h1 == coreId ? io_cache_coreResps_1_reqId_bits : io_cache_coreResps_0_reqId_bits; // @[Cat.scala 33:{92,92}]
  wire [1:0] _GEN_60 = 2'h2 == coreId ? io_cache_coreResps_2_reqId_bits : _GEN_59; // @[Cat.scala 33:{92,92}]
  wire [1:0] _GEN_61 = 2'h3 == coreId ? io_cache_coreResps_3_reqId_bits : _GEN_60; // @[Cat.scala 33:{92,92}]
  wire [2:0] _responseHead_T = {_GEN_57,_GEN_61}; // @[Cat.scala 33:92]
  wire [15:0] responseHead = {{13'd0}, _responseHead_T}; // @[CacheRequestController.scala 107:39 108:22]
  wire [7:0] _GEN_62 = _GEN_49 ? _GEN_53[7:0] : sendDataReg_0; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_63 = _GEN_49 ? _GEN_53[15:8] : sendDataReg_1; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_64 = _GEN_49 ? _GEN_53[23:16] : sendDataReg_2; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_65 = _GEN_49 ? _GEN_53[31:24] : sendDataReg_3; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_66 = _GEN_49 ? _GEN_53[39:32] : sendDataReg_4; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_67 = _GEN_49 ? _GEN_53[47:40] : sendDataReg_5; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_68 = _GEN_49 ? _GEN_53[55:48] : sendDataReg_6; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_69 = _GEN_49 ? _GEN_53[63:56] : sendDataReg_7; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_70 = _GEN_49 ? _GEN_53[71:64] : sendDataReg_8; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_71 = _GEN_49 ? _GEN_53[79:72] : sendDataReg_9; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_72 = _GEN_49 ? _GEN_53[87:80] : sendDataReg_10; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_73 = _GEN_49 ? _GEN_53[95:88] : sendDataReg_11; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_74 = _GEN_49 ? _GEN_53[103:96] : sendDataReg_12; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_75 = _GEN_49 ? _GEN_53[111:104] : sendDataReg_13; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_76 = _GEN_49 ? _GEN_53[119:112] : sendDataReg_14; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_77 = _GEN_49 ? _GEN_53[127:120] : sendDataReg_15; // @[CacheRequestController.scala 101:52 103:36 62:28]
  wire [7:0] _GEN_78 = _GEN_49 ? responseHead[7:0] : sendDataReg_16; // @[CacheRequestController.scala 101:52 110:53 62:28]
  wire [7:0] _GEN_79 = _GEN_49 ? responseHead[15:8] : sendDataReg_17; // @[CacheRequestController.scala 101:52 110:53 62:28]
  wire [1:0] _GEN_80 = _GEN_49 ? 2'h3 : stateReg; // @[CacheRequestController.scala 101:52 113:18 60:25]
  wire [4:0] _sendDataCntReg_T_1 = sendDataCntReg + 5'h1; // @[CacheRequestController.scala 120:42]
  wire [4:0] _GEN_81 = uart_io__txChannel_ready ? _sendDataCntReg_T_1 : sendDataCntReg; // @[CacheRequestController.scala 119:37 120:24 64:31]
  wire [1:0] _GEN_82 = sendDataCntReg == 5'h12 ? 2'h0 : stateReg; // @[CacheRequestController.scala 123:49 124:18 60:25]
  wire [4:0] _GEN_83 = sendDataCntReg == 5'h12 ? 5'h0 : _GEN_81; // @[CacheRequestController.scala 123:49 125:24]
  wire [4:0] _GEN_85 = 2'h3 == stateReg ? _GEN_83 : sendDataCntReg; // @[CacheRequestController.scala 80:20 64:31]
  wire [1:0] _GEN_86 = 2'h3 == stateReg ? _GEN_82 : stateReg; // @[CacheRequestController.scala 80:20 60:25]
  wire  _GEN_107 = 2'h2 == stateReg ? 1'h0 : 2'h3 == stateReg; // @[CacheRequestController.scala 80:20 66:28]
  wire  _GEN_130 = 2'h1 == stateReg ? 1'h0 : _GEN_107; // @[CacheRequestController.scala 80:20 66:28]
  wire  reqIdValid = rxReady ? 1'h0 : 2'h1 == stateReg; // @[CacheRequestController.scala 80:20 69:31]
  wire [7:0] _GEN_177 = 5'h1 == sendDataCntReg ? sendDataReg_1 : sendDataReg_0; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_178 = 5'h2 == sendDataCntReg ? sendDataReg_2 : _GEN_177; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_179 = 5'h3 == sendDataCntReg ? sendDataReg_3 : _GEN_178; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_180 = 5'h4 == sendDataCntReg ? sendDataReg_4 : _GEN_179; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_181 = 5'h5 == sendDataCntReg ? sendDataReg_5 : _GEN_180; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_182 = 5'h6 == sendDataCntReg ? sendDataReg_6 : _GEN_181; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_183 = 5'h7 == sendDataCntReg ? sendDataReg_7 : _GEN_182; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_184 = 5'h8 == sendDataCntReg ? sendDataReg_8 : _GEN_183; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_185 = 5'h9 == sendDataCntReg ? sendDataReg_9 : _GEN_184; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_186 = 5'ha == sendDataCntReg ? sendDataReg_10 : _GEN_185; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_187 = 5'hb == sendDataCntReg ? sendDataReg_11 : _GEN_186; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_188 = 5'hc == sendDataCntReg ? sendDataReg_12 : _GEN_187; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_189 = 5'hd == sendDataCntReg ? sendDataReg_13 : _GEN_188; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_190 = 5'he == sendDataCntReg ? sendDataReg_14 : _GEN_189; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_191 = 5'hf == sendDataCntReg ? sendDataReg_15 : _GEN_190; // @[CacheRequestController.scala 140:{10,10}]
  wire [7:0] _GEN_192 = 5'h10 == sendDataCntReg ? sendDataReg_16 : _GEN_191; // @[CacheRequestController.scala 140:{10,10}]
  Uart uart ( // @[CacheRequestController.scala 57:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io__rxd(uart_io__rxd),
    .io__txd(uart_io__txd),
    .io__rxChannel_ready(uart_io__rxChannel_ready),
    .io__rxChannel_valid(uart_io__rxChannel_valid),
    .io__rxChannel_bits(uart_io__rxChannel_bits),
    .io__txChannel_ready(uart_io__txChannel_ready),
    .io__txChannel_valid(uart_io__txChannel_valid),
    .io__txChannel_bits(uart_io__txChannel_bits)
  );
  assign io_txd = uart_io__txd; // @[CacheRequestController.scala 146:10]
  assign io_cache_coreReqs_0_reqId_valid = coreId == 2'h0 & reqIdValid; // @[CacheRequestController.scala 131:50]
  assign io_cache_coreReqs_0_reqId_bits = cmdAsUint[146:145]; // @[CacheRequestController.scala 75:24]
  assign io_cache_coreReqs_0_addr = cmdAsUint[142:128]; // @[CacheRequestController.scala 77:23]
  assign io_cache_coreReqs_0_rw = rw[0]; // @[CacheRequestController.scala 133:35]
  assign io_cache_coreReqs_0_wData = cmdAsUint[127:0]; // @[CacheRequestController.scala 78:24]
  assign io_cache_coreReqs_1_reqId_valid = coreId == 2'h1 & reqIdValid; // @[CacheRequestController.scala 131:50]
  assign io_cache_coreReqs_1_reqId_bits = cmdAsUint[146:145]; // @[CacheRequestController.scala 75:24]
  assign io_cache_coreReqs_1_addr = cmdAsUint[142:128]; // @[CacheRequestController.scala 77:23]
  assign io_cache_coreReqs_1_rw = rw[0]; // @[CacheRequestController.scala 133:35]
  assign io_cache_coreReqs_1_wData = cmdAsUint[127:0]; // @[CacheRequestController.scala 78:24]
  assign io_cache_coreReqs_2_reqId_valid = coreId == 2'h2 & reqIdValid; // @[CacheRequestController.scala 131:50]
  assign io_cache_coreReqs_2_reqId_bits = cmdAsUint[146:145]; // @[CacheRequestController.scala 75:24]
  assign io_cache_coreReqs_2_addr = cmdAsUint[142:128]; // @[CacheRequestController.scala 77:23]
  assign io_cache_coreReqs_2_rw = rw[0]; // @[CacheRequestController.scala 133:35]
  assign io_cache_coreReqs_2_wData = cmdAsUint[127:0]; // @[CacheRequestController.scala 78:24]
  assign io_cache_coreReqs_3_reqId_valid = coreId == 2'h3 & reqIdValid; // @[CacheRequestController.scala 131:50]
  assign io_cache_coreReqs_3_reqId_bits = cmdAsUint[146:145]; // @[CacheRequestController.scala 75:24]
  assign io_cache_coreReqs_3_addr = cmdAsUint[142:128]; // @[CacheRequestController.scala 77:23]
  assign io_cache_coreReqs_3_rw = rw[0]; // @[CacheRequestController.scala 133:35]
  assign io_cache_coreReqs_3_wData = cmdAsUint[127:0]; // @[CacheRequestController.scala 78:24]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io__rxd = io_rxd; // @[CacheRequestController.scala 147:15]
  assign uart_io__rxChannel_ready = 2'h0 == stateReg; // @[CacheRequestController.scala 80:20]
  assign uart_io__txChannel_valid = rxReady ? 1'h0 : _GEN_130; // @[CacheRequestController.scala 80:20 66:28]
  assign uart_io__txChannel_bits = 5'h11 == sendDataCntReg ? sendDataReg_17 : _GEN_192; // @[CacheRequestController.scala 140:{10,10}]
  always @(posedge clock) begin
    if (reset) begin // @[CacheRequestController.scala 60:25]
      stateReg <= 2'h0; // @[CacheRequestController.scala 60:25]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (cmdRcvCntReg == 5'h13) begin // @[CacheRequestController.scala 88:42]
        stateReg <= 2'h1; // @[CacheRequestController.scala 89:18]
      end
    end else if (2'h1 == stateReg) begin // @[CacheRequestController.scala 80:20]
      if (_GEN_44) begin // @[CacheRequestController.scala 95:51]
        stateReg <= 2'h2; // @[CacheRequestController.scala 96:18]
      end
    end else if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
      stateReg <= _GEN_80;
    end else begin
      stateReg <= _GEN_86;
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_0 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h0 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_0 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_1 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h1 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_1 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_2 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h2 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_2 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_3 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h3 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_3 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_4 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h4 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_4 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_5 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h5 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_5 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_6 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h6 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_6 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_7 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h7 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_7 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_8 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h8 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_8 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_9 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h9 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_9 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_10 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'ha == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_10 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_11 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'hb == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_11 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_12 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'hc == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_12 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_13 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'hd == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_13 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_14 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'he == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_14 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_15 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'hf == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_15 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_16 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h10 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_16 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_17 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h11 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_17 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 61:23]
      cmdReg_18 <= 8'h0; // @[CacheRequestController.scala 61:23]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        if (5'h12 == cmdRcvCntReg) begin // @[CacheRequestController.scala 85:30]
          cmdReg_18 <= _cmdReg_cmdRcvCntReg; // @[CacheRequestController.scala 85:30]
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_0 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_0 <= _GEN_62;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_1 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_1 <= _GEN_63;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_2 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_2 <= _GEN_64;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_3 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_3 <= _GEN_65;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_4 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_4 <= _GEN_66;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_5 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_5 <= _GEN_67;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_6 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_6 <= _GEN_68;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_7 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_7 <= _GEN_69;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_8 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_8 <= _GEN_70;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_9 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_9 <= _GEN_71;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_10 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_10 <= _GEN_72;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_11 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_11 <= _GEN_73;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_12 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_12 <= _GEN_74;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_13 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_13 <= _GEN_75;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_14 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_14 <= _GEN_76;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_15 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_15 <= _GEN_77;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_16 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_16 <= _GEN_78;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 62:28]
      sendDataReg_17 <= 8'h0; // @[CacheRequestController.scala 62:28]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (2'h2 == stateReg) begin // @[CacheRequestController.scala 80:20]
          sendDataReg_17 <= _GEN_79;
        end
      end
    end
    if (reset) begin // @[CacheRequestController.scala 63:29]
      cmdRcvCntReg <= 5'h0; // @[CacheRequestController.scala 63:29]
    end else if (rxReady) begin // @[CacheRequestController.scala 80:20]
      if (cmdRcvCntReg == 5'h13) begin // @[CacheRequestController.scala 88:42]
        cmdRcvCntReg <= 5'h0; // @[CacheRequestController.scala 90:22]
      end else if (uart_io__rxChannel_valid) begin // @[CacheRequestController.scala 83:37]
        cmdRcvCntReg <= _cmdRcvCntReg_T_1; // @[CacheRequestController.scala 84:22]
      end
    end
    if (reset) begin // @[CacheRequestController.scala 64:31]
      sendDataCntReg <= 5'h0; // @[CacheRequestController.scala 64:31]
    end else if (!(rxReady)) begin // @[CacheRequestController.scala 80:20]
      if (!(2'h1 == stateReg)) begin // @[CacheRequestController.scala 80:20]
        if (!(2'h2 == stateReg)) begin // @[CacheRequestController.scala 80:20]
          sendDataCntReg <= _GEN_85;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cmdReg_0 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  cmdReg_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  cmdReg_2 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  cmdReg_3 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  cmdReg_4 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  cmdReg_5 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  cmdReg_6 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  cmdReg_7 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  cmdReg_8 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  cmdReg_9 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  cmdReg_10 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  cmdReg_11 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  cmdReg_12 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  cmdReg_13 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  cmdReg_14 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  cmdReg_15 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  cmdReg_16 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  cmdReg_17 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  cmdReg_18 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  sendDataReg_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  sendDataReg_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  sendDataReg_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  sendDataReg_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  sendDataReg_4 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  sendDataReg_5 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  sendDataReg_6 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  sendDataReg_7 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  sendDataReg_8 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  sendDataReg_9 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  sendDataReg_10 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  sendDataReg_11 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  sendDataReg_12 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  sendDataReg_13 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  sendDataReg_14 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  sendDataReg_15 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  sendDataReg_16 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  sendDataReg_17 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  cmdRcvCntReg = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  sendDataCntReg = _RAND_39[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg  memReg_0; // @[RegFifo.scala 24:19]
  reg  memReg_1; // @[RegFifo.scala 24:19]
  reg  memReg_2; // @[RegFifo.scala 24:19]
  reg  memReg_3; // @[RegFifo.scala 24:19]
  reg  memReg_4; // @[RegFifo.scala 24:19]
  reg  memReg_5; // @[RegFifo.scala 24:19]
  reg  memReg_6; // @[RegFifo.scala 24:19]
  reg  memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire  _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire  _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire  _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire  _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire  _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_enq_ready = ~fullReg; // @[RegFifo.scala 82:19]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  always @(posedge clock) begin
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [1:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [1:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [1:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [1:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [1:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [1:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [1:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_enq_ready = ~fullReg; // @[RegFifo.scala 82:19]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  always @(posedge clock) begin
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo_3(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [127:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [127:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [127:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [127:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [127:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [127:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [127:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_enq_ready = ~fullReg; // @[RegFifo.scala 82:19]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  always @(posedge clock) begin
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  memReg_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  memReg_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  memReg_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  memReg_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  memReg_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  memReg_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  memReg_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  memReg_7 = _RAND_7[127:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo_4(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits,
  output [2:0] memReg_0_0,
  output [2:0] memReg_0_1,
  output [2:0] memReg_0_2,
  output [2:0] memReg_0_3,
  output [2:0] memReg_0_4,
  output [2:0] memReg_0_5,
  output [2:0] memReg_0_6,
  output [2:0] memReg_0_7,
  output [2:0] readPtr_0,
  output [2:0] writePtr_0,
  output       incrWrite_1,
  output       incrRead_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [2:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  doWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = doWrite; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [2:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [2:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [2:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [2:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [2:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [2:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_enq_ready = ~fullReg; // @[RegFifo.scala 82:19]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  assign memReg_0_0 = memReg_0;
  assign memReg_0_1 = memReg_1;
  assign memReg_0_2 = memReg_2;
  assign memReg_0_3 = memReg_3;
  assign memReg_0_4 = memReg_4;
  assign memReg_0_5 = memReg_5;
  assign memReg_0_6 = memReg_6;
  assign memReg_0_7 = memReg_7;
  assign readPtr_0 = readPtr;
  assign writePtr_0 = writePtr;
  assign incrWrite_1 = incrWrite;
  assign incrRead_0 = incrRead;
  always @(posedge clock) begin
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_3 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_5 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_6 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_7 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MshrQueue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits,
  output [2:0] io_regOut_0,
  output [2:0] io_regOut_1,
  output [2:0] io_regOut_2,
  output [2:0] io_regOut_3,
  output [2:0] io_regOut_4,
  output [2:0] io_regOut_5,
  output [2:0] io_regOut_6,
  output [2:0] io_regOut_7,
  output       io_validRegs_0,
  output       io_validRegs_1,
  output       io_validRegs_2,
  output       io_validRegs_3,
  output       io_validRegs_4,
  output       io_validRegs_5,
  output       io_validRegs_6,
  output       io_validRegs_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  fifo_clock; // @[MissFifo.scala 27:20]
  wire  fifo_reset; // @[MissFifo.scala 27:20]
  wire  fifo_io_enq_ready; // @[MissFifo.scala 27:20]
  wire  fifo_io_enq_valid; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_io_enq_bits; // @[MissFifo.scala 27:20]
  wire  fifo_io_deq_ready; // @[MissFifo.scala 27:20]
  wire  fifo_io_deq_valid; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_io_deq_bits; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_0; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_1; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_2; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_3; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_4; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_5; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_6; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_memReg_0_7; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_readPtr_0; // @[MissFifo.scala 27:20]
  wire [2:0] fifo_writePtr_0; // @[MissFifo.scala 27:20]
  wire  fifo_incrWrite_1; // @[MissFifo.scala 27:20]
  wire  fifo_incrRead_0; // @[MissFifo.scala 27:20]
  reg  validRegs_0; // @[MissFifo.scala 29:26]
  reg  validRegs_1; // @[MissFifo.scala 29:26]
  reg  validRegs_2; // @[MissFifo.scala 29:26]
  reg  validRegs_3; // @[MissFifo.scala 29:26]
  reg  validRegs_4; // @[MissFifo.scala 29:26]
  reg  validRegs_5; // @[MissFifo.scala 29:26]
  reg  validRegs_6; // @[MissFifo.scala 29:26]
  reg  validRegs_7; // @[MissFifo.scala 29:26]
  wire [2:0] readPtr = fifo_readPtr_0;
  wire  _GEN_0 = 3'h0 == readPtr ? 1'h0 : validRegs_0; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_1 = 3'h1 == readPtr ? 1'h0 : validRegs_1; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_2 = 3'h2 == readPtr ? 1'h0 : validRegs_2; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_3 = 3'h3 == readPtr ? 1'h0 : validRegs_3; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_4 = 3'h4 == readPtr ? 1'h0 : validRegs_4; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_5 = 3'h5 == readPtr ? 1'h0 : validRegs_5; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_6 = 3'h6 == readPtr ? 1'h0 : validRegs_6; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  _GEN_7 = 3'h7 == readPtr ? 1'h0 : validRegs_7; // @[MissFifo.scala 43:{22,22} 29:26]
  wire  incrRead_0 = fifo_incrRead_0;
  wire  _GEN_8 = incrRead_0 ? _GEN_0 : validRegs_0; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_9 = incrRead_0 ? _GEN_1 : validRegs_1; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_10 = incrRead_0 ? _GEN_2 : validRegs_2; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_11 = incrRead_0 ? _GEN_3 : validRegs_3; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_12 = incrRead_0 ? _GEN_4 : validRegs_4; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_13 = incrRead_0 ? _GEN_5 : validRegs_5; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_14 = incrRead_0 ? _GEN_6 : validRegs_6; // @[MissFifo.scala 42:18 29:26]
  wire  _GEN_15 = incrRead_0 ? _GEN_7 : validRegs_7; // @[MissFifo.scala 42:18 29:26]
  wire [2:0] writePtr = fifo_writePtr_0;
  wire  _GEN_16 = 3'h0 == writePtr | _GEN_8; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_17 = 3'h1 == writePtr | _GEN_9; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_18 = 3'h2 == writePtr | _GEN_10; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_19 = 3'h3 == writePtr | _GEN_11; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_20 = 3'h4 == writePtr | _GEN_12; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_21 = 3'h5 == writePtr | _GEN_13; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_22 = 3'h6 == writePtr | _GEN_14; // @[MissFifo.scala 47:{22,22}]
  wire  _GEN_23 = 3'h7 == writePtr | _GEN_15; // @[MissFifo.scala 47:{22,22}]
  wire  incrWrite_1 = fifo_incrWrite_1;
  RegFifo_4 fifo ( // @[MissFifo.scala 27:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .memReg_0_0(fifo_memReg_0_0),
    .memReg_0_1(fifo_memReg_0_1),
    .memReg_0_2(fifo_memReg_0_2),
    .memReg_0_3(fifo_memReg_0_3),
    .memReg_0_4(fifo_memReg_0_4),
    .memReg_0_5(fifo_memReg_0_5),
    .memReg_0_6(fifo_memReg_0_6),
    .memReg_0_7(fifo_memReg_0_7),
    .readPtr_0(fifo_readPtr_0),
    .writePtr_0(fifo_writePtr_0),
    .incrWrite_1(fifo_incrWrite_1),
    .incrRead_0(fifo_incrRead_0)
  );
  assign io_enq_ready = fifo_io_enq_ready; // @[MissFifo.scala 53:10]
  assign io_deq_valid = fifo_io_deq_valid; // @[MissFifo.scala 52:10]
  assign io_deq_bits = fifo_io_deq_bits; // @[MissFifo.scala 52:10]
  assign io_regOut_0 = fifo_memReg_0_0; // @[MissFifo.scala 28:23]
  assign io_regOut_1 = fifo_memReg_0_1; // @[MissFifo.scala 28:23]
  assign io_regOut_2 = fifo_memReg_0_2; // @[MissFifo.scala 28:23]
  assign io_regOut_3 = fifo_memReg_0_3; // @[MissFifo.scala 28:23]
  assign io_regOut_4 = fifo_memReg_0_4; // @[MissFifo.scala 28:23]
  assign io_regOut_5 = fifo_memReg_0_5; // @[MissFifo.scala 28:23]
  assign io_regOut_6 = fifo_memReg_0_6; // @[MissFifo.scala 28:23]
  assign io_regOut_7 = fifo_memReg_0_7; // @[MissFifo.scala 28:23]
  assign io_validRegs_0 = validRegs_0; // @[MissFifo.scala 50:16]
  assign io_validRegs_1 = validRegs_1; // @[MissFifo.scala 50:16]
  assign io_validRegs_2 = validRegs_2; // @[MissFifo.scala 50:16]
  assign io_validRegs_3 = validRegs_3; // @[MissFifo.scala 50:16]
  assign io_validRegs_4 = validRegs_4; // @[MissFifo.scala 50:16]
  assign io_validRegs_5 = validRegs_5; // @[MissFifo.scala 50:16]
  assign io_validRegs_6 = validRegs_6; // @[MissFifo.scala 50:16]
  assign io_validRegs_7 = validRegs_7; // @[MissFifo.scala 50:16]
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_enq_valid = io_enq_valid; // @[MissFifo.scala 53:10]
  assign fifo_io_enq_bits = io_enq_bits; // @[MissFifo.scala 53:10]
  assign fifo_io_deq_ready = io_deq_ready; // @[MissFifo.scala 52:10]
  always @(posedge clock) begin
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_0 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_0 <= _GEN_16;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h0 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_0 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_1 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_1 <= _GEN_17;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h1 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_1 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_2 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_2 <= _GEN_18;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h2 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_2 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_3 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_3 <= _GEN_19;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h3 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_3 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_4 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_4 <= _GEN_20;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h4 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_4 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_5 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_5 <= _GEN_21;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h5 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_5 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_6 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_6 <= _GEN_22;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h6 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_6 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
    if (reset) begin // @[MissFifo.scala 29:26]
      validRegs_7 <= 1'h0; // @[MissFifo.scala 29:26]
    end else if (incrWrite_1) begin // @[MissFifo.scala 46:19]
      validRegs_7 <= _GEN_23;
    end else if (incrRead_0) begin // @[MissFifo.scala 42:18]
      if (3'h7 == readPtr) begin // @[MissFifo.scala 43:22]
        validRegs_7 <= 1'h0; // @[MissFifo.scala 43:22]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validRegs_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  validRegs_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  validRegs_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  validRegs_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  validRegs_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  validRegs_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  validRegs_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  validRegs_7 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo_5(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [3:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [3:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_enq_ready = ~fullReg; // @[RegFifo.scala 82:19]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  always @(posedge clock) begin
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo_6(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [4:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [4:0] io_deq_bits,
  output [4:0] memReg_1_0,
  output [4:0] memReg_1_1,
  output [4:0] memReg_1_2,
  output [4:0] memReg_1_3,
  output [4:0] memReg_1_4,
  output [4:0] memReg_1_5,
  output [4:0] memReg_1_6,
  output [4:0] memReg_1_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  doWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = doWrite; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [4:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_enq_ready = ~fullReg; // @[RegFifo.scala 82:19]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  assign memReg_1_0 = memReg_0;
  assign memReg_1_1 = memReg_1;
  assign memReg_1_2 = memReg_2;
  assign memReg_1_3 = memReg_3;
  assign memReg_1_4 = memReg_4;
  assign memReg_1_5 = memReg_5;
  assign memReg_1_6 = memReg_6;
  assign memReg_1_7 = memReg_7;
  always @(posedge clock) begin
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (doWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_4 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_5 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_6 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_7 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MshrQueue_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [4:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [4:0] io_deq_bits,
  output [4:0] io_regOut_0,
  output [4:0] io_regOut_1,
  output [4:0] io_regOut_2,
  output [4:0] io_regOut_3,
  output [4:0] io_regOut_4,
  output [4:0] io_regOut_5,
  output [4:0] io_regOut_6,
  output [4:0] io_regOut_7
);
  wire  fifo_clock; // @[MissFifo.scala 27:20]
  wire  fifo_reset; // @[MissFifo.scala 27:20]
  wire  fifo_io_enq_ready; // @[MissFifo.scala 27:20]
  wire  fifo_io_enq_valid; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_io_enq_bits; // @[MissFifo.scala 27:20]
  wire  fifo_io_deq_ready; // @[MissFifo.scala 27:20]
  wire  fifo_io_deq_valid; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_io_deq_bits; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_0; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_1; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_2; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_3; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_4; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_5; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_6; // @[MissFifo.scala 27:20]
  wire [4:0] fifo_memReg_1_7; // @[MissFifo.scala 27:20]
  RegFifo_6 fifo ( // @[MissFifo.scala 27:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .memReg_1_0(fifo_memReg_1_0),
    .memReg_1_1(fifo_memReg_1_1),
    .memReg_1_2(fifo_memReg_1_2),
    .memReg_1_3(fifo_memReg_1_3),
    .memReg_1_4(fifo_memReg_1_4),
    .memReg_1_5(fifo_memReg_1_5),
    .memReg_1_6(fifo_memReg_1_6),
    .memReg_1_7(fifo_memReg_1_7)
  );
  assign io_enq_ready = fifo_io_enq_ready; // @[MissFifo.scala 53:10]
  assign io_deq_valid = fifo_io_deq_valid; // @[MissFifo.scala 52:10]
  assign io_deq_bits = fifo_io_deq_bits; // @[MissFifo.scala 52:10]
  assign io_regOut_0 = fifo_memReg_1_0; // @[MissFifo.scala 28:23]
  assign io_regOut_1 = fifo_memReg_1_1; // @[MissFifo.scala 28:23]
  assign io_regOut_2 = fifo_memReg_1_2; // @[MissFifo.scala 28:23]
  assign io_regOut_3 = fifo_memReg_1_3; // @[MissFifo.scala 28:23]
  assign io_regOut_4 = fifo_memReg_1_4; // @[MissFifo.scala 28:23]
  assign io_regOut_5 = fifo_memReg_1_5; // @[MissFifo.scala 28:23]
  assign io_regOut_6 = fifo_memReg_1_6; // @[MissFifo.scala 28:23]
  assign io_regOut_7 = fifo_memReg_1_7; // @[MissFifo.scala 28:23]
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_enq_valid = io_enq_valid; // @[MissFifo.scala 53:10]
  assign fifo_io_enq_bits = io_enq_bits; // @[MissFifo.scala 53:10]
  assign fifo_io_deq_ready = io_deq_ready; // @[MissFifo.scala 52:10]
endmodule
module MissFifo(
  input          clock,
  input          reset,
  input          io_push,
  input          io_pushEntry_rw,
  input  [1:0]   io_pushEntry_reqId,
  input  [1:0]   io_pushEntry_coreId,
  input  [127:0] io_pushEntry_wData,
  input  [2:0]   io_pushEntry_replaceWay,
  input  [3:0]   io_pushEntry_tag,
  input  [4:0]   io_pushEntry_index,
  input  [1:0]   io_pushEntry_blockOffset,
  input          io_pop,
  output         io_popEntry_rw,
  output [1:0]   io_popEntry_reqId,
  output [1:0]   io_popEntry_coreId,
  output [127:0] io_popEntry_wData,
  output [2:0]   io_popEntry_replaceWay,
  output [3:0]   io_popEntry_tag,
  output [4:0]   io_popEntry_index,
  output [1:0]   io_popEntry_blockOffset,
  output [4:0]   io_currentIndexes_0,
  output [4:0]   io_currentIndexes_1,
  output [4:0]   io_currentIndexes_2,
  output [4:0]   io_currentIndexes_3,
  output [4:0]   io_currentIndexes_4,
  output [4:0]   io_currentIndexes_5,
  output [4:0]   io_currentIndexes_6,
  output [4:0]   io_currentIndexes_7,
  output [2:0]   io_currentWays_0,
  output [2:0]   io_currentWays_1,
  output [2:0]   io_currentWays_2,
  output [2:0]   io_currentWays_3,
  output [2:0]   io_currentWays_4,
  output [2:0]   io_currentWays_5,
  output [2:0]   io_currentWays_6,
  output [2:0]   io_currentWays_7,
  output         io_validMSHRs_0,
  output         io_validMSHRs_1,
  output         io_validMSHRs_2,
  output         io_validMSHRs_3,
  output         io_validMSHRs_4,
  output         io_validMSHRs_5,
  output         io_validMSHRs_6,
  output         io_validMSHRs_7,
  output         io_full,
  output         io_empty
);
  wire  rwQueue_clock; // @[MissFifo.scala 69:23]
  wire  rwQueue_reset; // @[MissFifo.scala 69:23]
  wire  rwQueue_io_enq_ready; // @[MissFifo.scala 69:23]
  wire  rwQueue_io_enq_valid; // @[MissFifo.scala 69:23]
  wire  rwQueue_io_enq_bits; // @[MissFifo.scala 69:23]
  wire  rwQueue_io_deq_ready; // @[MissFifo.scala 69:23]
  wire  rwQueue_io_deq_valid; // @[MissFifo.scala 69:23]
  wire  rwQueue_io_deq_bits; // @[MissFifo.scala 69:23]
  wire  reqIdQueue_clock; // @[MissFifo.scala 70:26]
  wire  reqIdQueue_reset; // @[MissFifo.scala 70:26]
  wire  reqIdQueue_io_enq_ready; // @[MissFifo.scala 70:26]
  wire  reqIdQueue_io_enq_valid; // @[MissFifo.scala 70:26]
  wire [1:0] reqIdQueue_io_enq_bits; // @[MissFifo.scala 70:26]
  wire  reqIdQueue_io_deq_ready; // @[MissFifo.scala 70:26]
  wire  reqIdQueue_io_deq_valid; // @[MissFifo.scala 70:26]
  wire [1:0] reqIdQueue_io_deq_bits; // @[MissFifo.scala 70:26]
  wire  coreIdQueue_clock; // @[MissFifo.scala 71:27]
  wire  coreIdQueue_reset; // @[MissFifo.scala 71:27]
  wire  coreIdQueue_io_enq_ready; // @[MissFifo.scala 71:27]
  wire  coreIdQueue_io_enq_valid; // @[MissFifo.scala 71:27]
  wire [1:0] coreIdQueue_io_enq_bits; // @[MissFifo.scala 71:27]
  wire  coreIdQueue_io_deq_ready; // @[MissFifo.scala 71:27]
  wire  coreIdQueue_io_deq_valid; // @[MissFifo.scala 71:27]
  wire [1:0] coreIdQueue_io_deq_bits; // @[MissFifo.scala 71:27]
  wire  wDataQueue_clock; // @[MissFifo.scala 72:26]
  wire  wDataQueue_reset; // @[MissFifo.scala 72:26]
  wire  wDataQueue_io_enq_ready; // @[MissFifo.scala 72:26]
  wire  wDataQueue_io_enq_valid; // @[MissFifo.scala 72:26]
  wire [127:0] wDataQueue_io_enq_bits; // @[MissFifo.scala 72:26]
  wire  wDataQueue_io_deq_ready; // @[MissFifo.scala 72:26]
  wire  wDataQueue_io_deq_valid; // @[MissFifo.scala 72:26]
  wire [127:0] wDataQueue_io_deq_bits; // @[MissFifo.scala 72:26]
  wire  wayQueue_clock; // @[MissFifo.scala 73:24]
  wire  wayQueue_reset; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_enq_ready; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_enq_valid; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_enq_bits; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_deq_ready; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_deq_valid; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_deq_bits; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_0; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_1; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_2; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_3; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_4; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_5; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_6; // @[MissFifo.scala 73:24]
  wire [2:0] wayQueue_io_regOut_7; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_0; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_1; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_2; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_3; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_4; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_5; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_6; // @[MissFifo.scala 73:24]
  wire  wayQueue_io_validRegs_7; // @[MissFifo.scala 73:24]
  wire  tagQueue_clock; // @[MissFifo.scala 74:24]
  wire  tagQueue_reset; // @[MissFifo.scala 74:24]
  wire  tagQueue_io_enq_ready; // @[MissFifo.scala 74:24]
  wire  tagQueue_io_enq_valid; // @[MissFifo.scala 74:24]
  wire [3:0] tagQueue_io_enq_bits; // @[MissFifo.scala 74:24]
  wire  tagQueue_io_deq_ready; // @[MissFifo.scala 74:24]
  wire  tagQueue_io_deq_valid; // @[MissFifo.scala 74:24]
  wire [3:0] tagQueue_io_deq_bits; // @[MissFifo.scala 74:24]
  wire  idxQueue_clock; // @[MissFifo.scala 75:24]
  wire  idxQueue_reset; // @[MissFifo.scala 75:24]
  wire  idxQueue_io_enq_ready; // @[MissFifo.scala 75:24]
  wire  idxQueue_io_enq_valid; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_enq_bits; // @[MissFifo.scala 75:24]
  wire  idxQueue_io_deq_ready; // @[MissFifo.scala 75:24]
  wire  idxQueue_io_deq_valid; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_deq_bits; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_0; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_1; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_2; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_3; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_4; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_5; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_6; // @[MissFifo.scala 75:24]
  wire [4:0] idxQueue_io_regOut_7; // @[MissFifo.scala 75:24]
  wire  blockOffQueue_clock; // @[MissFifo.scala 76:29]
  wire  blockOffQueue_reset; // @[MissFifo.scala 76:29]
  wire  blockOffQueue_io_enq_ready; // @[MissFifo.scala 76:29]
  wire  blockOffQueue_io_enq_valid; // @[MissFifo.scala 76:29]
  wire [1:0] blockOffQueue_io_enq_bits; // @[MissFifo.scala 76:29]
  wire  blockOffQueue_io_deq_ready; // @[MissFifo.scala 76:29]
  wire  blockOffQueue_io_deq_valid; // @[MissFifo.scala 76:29]
  wire [1:0] blockOffQueue_io_deq_bits; // @[MissFifo.scala 76:29]
  wire  _full_T_1 = ~reqIdQueue_io_enq_ready; // @[MissFifo.scala 79:14]
  wire  _full_T_2 = ~rwQueue_io_enq_ready | _full_T_1; // @[MissFifo.scala 78:36]
  wire  _full_T_3 = ~coreIdQueue_io_enq_ready; // @[MissFifo.scala 80:14]
  wire  _full_T_4 = _full_T_2 | _full_T_3; // @[MissFifo.scala 79:39]
  wire  _full_T_5 = ~wDataQueue_io_enq_ready; // @[MissFifo.scala 81:14]
  wire  _full_T_6 = _full_T_4 | _full_T_5; // @[MissFifo.scala 80:40]
  wire  _full_T_7 = ~wayQueue_io_enq_ready; // @[MissFifo.scala 82:14]
  wire  _full_T_8 = _full_T_6 | _full_T_7; // @[MissFifo.scala 81:39]
  wire  _full_T_9 = ~tagQueue_io_enq_ready; // @[MissFifo.scala 83:14]
  wire  _full_T_10 = _full_T_8 | _full_T_9; // @[MissFifo.scala 82:37]
  wire  _full_T_11 = ~idxQueue_io_enq_ready; // @[MissFifo.scala 84:14]
  wire  _full_T_12 = _full_T_10 | _full_T_11; // @[MissFifo.scala 83:37]
  wire  _full_T_13 = ~blockOffQueue_io_enq_ready; // @[MissFifo.scala 85:14]
  wire  _empty_T_1 = ~reqIdQueue_io_deq_valid; // @[MissFifo.scala 88:15]
  wire  _empty_T_2 = ~rwQueue_io_deq_valid | _empty_T_1; // @[MissFifo.scala 87:37]
  wire  _empty_T_3 = ~coreIdQueue_io_deq_valid; // @[MissFifo.scala 89:15]
  wire  _empty_T_4 = _empty_T_2 | _empty_T_3; // @[MissFifo.scala 88:40]
  wire  _empty_T_5 = ~wDataQueue_io_deq_valid; // @[MissFifo.scala 90:15]
  wire  _empty_T_6 = _empty_T_4 | _empty_T_5; // @[MissFifo.scala 89:41]
  wire  _empty_T_7 = ~wayQueue_io_deq_valid; // @[MissFifo.scala 91:15]
  wire  _empty_T_8 = _empty_T_6 | _empty_T_7; // @[MissFifo.scala 90:40]
  wire  _empty_T_9 = ~tagQueue_io_deq_valid; // @[MissFifo.scala 92:15]
  wire  _empty_T_10 = _empty_T_8 | _empty_T_9; // @[MissFifo.scala 91:38]
  wire  _empty_T_11 = ~idxQueue_io_deq_valid; // @[MissFifo.scala 93:15]
  wire  _empty_T_12 = _empty_T_10 | _empty_T_11; // @[MissFifo.scala 92:38]
  wire  _empty_T_13 = ~blockOffQueue_io_deq_valid; // @[MissFifo.scala 94:15]
  RegFifo rwQueue ( // @[MissFifo.scala 69:23]
    .clock(rwQueue_clock),
    .reset(rwQueue_reset),
    .io_enq_ready(rwQueue_io_enq_ready),
    .io_enq_valid(rwQueue_io_enq_valid),
    .io_enq_bits(rwQueue_io_enq_bits),
    .io_deq_ready(rwQueue_io_deq_ready),
    .io_deq_valid(rwQueue_io_deq_valid),
    .io_deq_bits(rwQueue_io_deq_bits)
  );
  RegFifo_1 reqIdQueue ( // @[MissFifo.scala 70:26]
    .clock(reqIdQueue_clock),
    .reset(reqIdQueue_reset),
    .io_enq_ready(reqIdQueue_io_enq_ready),
    .io_enq_valid(reqIdQueue_io_enq_valid),
    .io_enq_bits(reqIdQueue_io_enq_bits),
    .io_deq_ready(reqIdQueue_io_deq_ready),
    .io_deq_valid(reqIdQueue_io_deq_valid),
    .io_deq_bits(reqIdQueue_io_deq_bits)
  );
  RegFifo_1 coreIdQueue ( // @[MissFifo.scala 71:27]
    .clock(coreIdQueue_clock),
    .reset(coreIdQueue_reset),
    .io_enq_ready(coreIdQueue_io_enq_ready),
    .io_enq_valid(coreIdQueue_io_enq_valid),
    .io_enq_bits(coreIdQueue_io_enq_bits),
    .io_deq_ready(coreIdQueue_io_deq_ready),
    .io_deq_valid(coreIdQueue_io_deq_valid),
    .io_deq_bits(coreIdQueue_io_deq_bits)
  );
  RegFifo_3 wDataQueue ( // @[MissFifo.scala 72:26]
    .clock(wDataQueue_clock),
    .reset(wDataQueue_reset),
    .io_enq_ready(wDataQueue_io_enq_ready),
    .io_enq_valid(wDataQueue_io_enq_valid),
    .io_enq_bits(wDataQueue_io_enq_bits),
    .io_deq_ready(wDataQueue_io_deq_ready),
    .io_deq_valid(wDataQueue_io_deq_valid),
    .io_deq_bits(wDataQueue_io_deq_bits)
  );
  MshrQueue wayQueue ( // @[MissFifo.scala 73:24]
    .clock(wayQueue_clock),
    .reset(wayQueue_reset),
    .io_enq_ready(wayQueue_io_enq_ready),
    .io_enq_valid(wayQueue_io_enq_valid),
    .io_enq_bits(wayQueue_io_enq_bits),
    .io_deq_ready(wayQueue_io_deq_ready),
    .io_deq_valid(wayQueue_io_deq_valid),
    .io_deq_bits(wayQueue_io_deq_bits),
    .io_regOut_0(wayQueue_io_regOut_0),
    .io_regOut_1(wayQueue_io_regOut_1),
    .io_regOut_2(wayQueue_io_regOut_2),
    .io_regOut_3(wayQueue_io_regOut_3),
    .io_regOut_4(wayQueue_io_regOut_4),
    .io_regOut_5(wayQueue_io_regOut_5),
    .io_regOut_6(wayQueue_io_regOut_6),
    .io_regOut_7(wayQueue_io_regOut_7),
    .io_validRegs_0(wayQueue_io_validRegs_0),
    .io_validRegs_1(wayQueue_io_validRegs_1),
    .io_validRegs_2(wayQueue_io_validRegs_2),
    .io_validRegs_3(wayQueue_io_validRegs_3),
    .io_validRegs_4(wayQueue_io_validRegs_4),
    .io_validRegs_5(wayQueue_io_validRegs_5),
    .io_validRegs_6(wayQueue_io_validRegs_6),
    .io_validRegs_7(wayQueue_io_validRegs_7)
  );
  RegFifo_5 tagQueue ( // @[MissFifo.scala 74:24]
    .clock(tagQueue_clock),
    .reset(tagQueue_reset),
    .io_enq_ready(tagQueue_io_enq_ready),
    .io_enq_valid(tagQueue_io_enq_valid),
    .io_enq_bits(tagQueue_io_enq_bits),
    .io_deq_ready(tagQueue_io_deq_ready),
    .io_deq_valid(tagQueue_io_deq_valid),
    .io_deq_bits(tagQueue_io_deq_bits)
  );
  MshrQueue_1 idxQueue ( // @[MissFifo.scala 75:24]
    .clock(idxQueue_clock),
    .reset(idxQueue_reset),
    .io_enq_ready(idxQueue_io_enq_ready),
    .io_enq_valid(idxQueue_io_enq_valid),
    .io_enq_bits(idxQueue_io_enq_bits),
    .io_deq_ready(idxQueue_io_deq_ready),
    .io_deq_valid(idxQueue_io_deq_valid),
    .io_deq_bits(idxQueue_io_deq_bits),
    .io_regOut_0(idxQueue_io_regOut_0),
    .io_regOut_1(idxQueue_io_regOut_1),
    .io_regOut_2(idxQueue_io_regOut_2),
    .io_regOut_3(idxQueue_io_regOut_3),
    .io_regOut_4(idxQueue_io_regOut_4),
    .io_regOut_5(idxQueue_io_regOut_5),
    .io_regOut_6(idxQueue_io_regOut_6),
    .io_regOut_7(idxQueue_io_regOut_7)
  );
  RegFifo_1 blockOffQueue ( // @[MissFifo.scala 76:29]
    .clock(blockOffQueue_clock),
    .reset(blockOffQueue_reset),
    .io_enq_ready(blockOffQueue_io_enq_ready),
    .io_enq_valid(blockOffQueue_io_enq_valid),
    .io_enq_bits(blockOffQueue_io_enq_bits),
    .io_deq_ready(blockOffQueue_io_deq_ready),
    .io_deq_valid(blockOffQueue_io_deq_valid),
    .io_deq_bits(blockOffQueue_io_deq_bits)
  );
  assign io_popEntry_rw = rwQueue_io_deq_bits; // @[MissFifo.scala 133:18]
  assign io_popEntry_reqId = reqIdQueue_io_deq_bits; // @[MissFifo.scala 134:21]
  assign io_popEntry_coreId = coreIdQueue_io_deq_bits; // @[MissFifo.scala 135:22]
  assign io_popEntry_wData = wDataQueue_io_deq_bits; // @[MissFifo.scala 136:21]
  assign io_popEntry_replaceWay = wayQueue_io_deq_bits; // @[MissFifo.scala 137:26]
  assign io_popEntry_tag = tagQueue_io_deq_bits; // @[MissFifo.scala 138:19]
  assign io_popEntry_index = idxQueue_io_deq_bits; // @[MissFifo.scala 139:21]
  assign io_popEntry_blockOffset = blockOffQueue_io_deq_bits; // @[MissFifo.scala 140:27]
  assign io_currentIndexes_0 = idxQueue_io_regOut_0; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_1 = idxQueue_io_regOut_1; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_2 = idxQueue_io_regOut_2; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_3 = idxQueue_io_regOut_3; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_4 = idxQueue_io_regOut_4; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_5 = idxQueue_io_regOut_5; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_6 = idxQueue_io_regOut_6; // @[MissFifo.scala 126:26]
  assign io_currentIndexes_7 = idxQueue_io_regOut_7; // @[MissFifo.scala 126:26]
  assign io_currentWays_0 = wayQueue_io_regOut_0; // @[MissFifo.scala 125:23]
  assign io_currentWays_1 = wayQueue_io_regOut_1; // @[MissFifo.scala 125:23]
  assign io_currentWays_2 = wayQueue_io_regOut_2; // @[MissFifo.scala 125:23]
  assign io_currentWays_3 = wayQueue_io_regOut_3; // @[MissFifo.scala 125:23]
  assign io_currentWays_4 = wayQueue_io_regOut_4; // @[MissFifo.scala 125:23]
  assign io_currentWays_5 = wayQueue_io_regOut_5; // @[MissFifo.scala 125:23]
  assign io_currentWays_6 = wayQueue_io_regOut_6; // @[MissFifo.scala 125:23]
  assign io_currentWays_7 = wayQueue_io_regOut_7; // @[MissFifo.scala 125:23]
  assign io_validMSHRs_0 = wayQueue_io_validRegs_0; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_1 = wayQueue_io_validRegs_1; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_2 = wayQueue_io_validRegs_2; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_3 = wayQueue_io_validRegs_3; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_4 = wayQueue_io_validRegs_4; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_5 = wayQueue_io_validRegs_5; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_6 = wayQueue_io_validRegs_6; // @[MissFifo.scala 132:17]
  assign io_validMSHRs_7 = wayQueue_io_validRegs_7; // @[MissFifo.scala 132:17]
  assign io_full = _full_T_12 | _full_T_13; // @[MissFifo.scala 84:37]
  assign io_empty = _empty_T_12 | _empty_T_13; // @[MissFifo.scala 93:38]
  assign rwQueue_clock = clock;
  assign rwQueue_reset = reset;
  assign rwQueue_io_enq_valid = io_push; // @[MissFifo.scala 97:24]
  assign rwQueue_io_enq_bits = io_pushEntry_rw; // @[MissFifo.scala 98:23]
  assign rwQueue_io_deq_ready = io_pop; // @[MissFifo.scala 115:24]
  assign reqIdQueue_clock = clock;
  assign reqIdQueue_reset = reset;
  assign reqIdQueue_io_enq_valid = io_push; // @[MissFifo.scala 99:27]
  assign reqIdQueue_io_enq_bits = io_pushEntry_reqId; // @[MissFifo.scala 100:26]
  assign reqIdQueue_io_deq_ready = io_pop; // @[MissFifo.scala 116:27]
  assign coreIdQueue_clock = clock;
  assign coreIdQueue_reset = reset;
  assign coreIdQueue_io_enq_valid = io_push; // @[MissFifo.scala 101:28]
  assign coreIdQueue_io_enq_bits = io_pushEntry_coreId; // @[MissFifo.scala 102:27]
  assign coreIdQueue_io_deq_ready = io_pop; // @[MissFifo.scala 117:28]
  assign wDataQueue_clock = clock;
  assign wDataQueue_reset = reset;
  assign wDataQueue_io_enq_valid = io_push; // @[MissFifo.scala 103:27]
  assign wDataQueue_io_enq_bits = io_pushEntry_wData; // @[MissFifo.scala 104:26]
  assign wDataQueue_io_deq_ready = io_pop; // @[MissFifo.scala 118:27]
  assign wayQueue_clock = clock;
  assign wayQueue_reset = reset;
  assign wayQueue_io_enq_valid = io_push; // @[MissFifo.scala 105:25]
  assign wayQueue_io_enq_bits = io_pushEntry_replaceWay; // @[MissFifo.scala 106:24]
  assign wayQueue_io_deq_ready = io_pop; // @[MissFifo.scala 119:25]
  assign tagQueue_clock = clock;
  assign tagQueue_reset = reset;
  assign tagQueue_io_enq_valid = io_push; // @[MissFifo.scala 107:25]
  assign tagQueue_io_enq_bits = io_pushEntry_tag; // @[MissFifo.scala 108:24]
  assign tagQueue_io_deq_ready = io_pop; // @[MissFifo.scala 120:25]
  assign idxQueue_clock = clock;
  assign idxQueue_reset = reset;
  assign idxQueue_io_enq_valid = io_push; // @[MissFifo.scala 109:25]
  assign idxQueue_io_enq_bits = io_pushEntry_index; // @[MissFifo.scala 110:24]
  assign idxQueue_io_deq_ready = io_pop; // @[MissFifo.scala 121:25]
  assign blockOffQueue_clock = clock;
  assign blockOffQueue_reset = reset;
  assign blockOffQueue_io_enq_valid = io_push; // @[MissFifo.scala 111:30]
  assign blockOffQueue_io_enq_bits = io_pushEntry_blockOffset; // @[MissFifo.scala 112:29]
  assign blockOffQueue_io_deq_ready = io_pop; // @[MissFifo.scala 122:30]
endmodule
module UpdateUnit(
  input          io_readStage_valid,
  input  [1:0]   io_readStage_reqId,
  input  [1:0]   io_readStage_coreId,
  input          io_readStage_rw,
  input  [127:0] io_readStage_wData,
  input  [2:0]   io_readStage_wWay,
  input  [3:0]   io_readStage_tag,
  input  [4:0]   io_readStage_index,
  input  [1:0]   io_readStage_blockOffset,
  input  [127:0] io_readStage_memReadData_0,
  input  [127:0] io_readStage_memReadData_1,
  input  [127:0] io_readStage_memReadData_2,
  input  [127:0] io_readStage_memReadData_3,
  input          io_memoryInterface_valid,
  input  [1:0]   io_memoryInterface_reqId,
  input  [1:0]   io_memoryInterface_coreId,
  input          io_memoryInterface_rw,
  input  [127:0] io_memoryInterface_wData,
  input  [2:0]   io_memoryInterface_wWay,
  input          io_memoryInterface_responseStatus,
  input  [3:0]   io_memoryInterface_tag,
  input  [4:0]   io_memoryInterface_index,
  input  [1:0]   io_memoryInterface_blockOffset,
  input  [127:0] io_memoryInterface_memReadData_0,
  input  [127:0] io_memoryInterface_memReadData_1,
  input  [127:0] io_memoryInterface_memReadData_2,
  input  [127:0] io_memoryInterface_memReadData_3,
  output [3:0]   io_cacheUpdateControl_tag,
  output [2:0]   io_cacheUpdateControl_index,
  output [1:0]   io_cacheUpdateControl_coreId,
  output [2:0]   io_cacheUpdateControl_way,
  output         io_cacheUpdateControl_refill,
  output         io_cacheUpdateControl_update,
  output         io_cacheUpdateControl_stall,
  output [127:0] io_cacheUpdateControl_memWriteData_0,
  output [127:0] io_cacheUpdateControl_memWriteData_1,
  output [127:0] io_cacheUpdateControl_memWriteData_2,
  output [127:0] io_cacheUpdateControl_memWriteData_3,
  output         io_cacheUpdateControl_wrEn,
  output         io_coreResp_reqId_valid,
  output [1:0]   io_coreResp_reqId_bits,
  output [127:0] io_coreResp_rData,
  output         io_coreResp_responseStatus
);
  wire [127:0] _cacheWriteData_0_T_1 = io_memoryInterface_blockOffset == 2'h0 ? io_memoryInterface_wData :
    io_memoryInterface_memReadData_0; // @[UpdateUnit.scala 68:33]
  wire [127:0] _cacheWriteData_1_T_1 = io_memoryInterface_blockOffset == 2'h1 ? io_memoryInterface_wData :
    io_memoryInterface_memReadData_1; // @[UpdateUnit.scala 68:33]
  wire [127:0] _cacheWriteData_2_T_1 = io_memoryInterface_blockOffset == 2'h2 ? io_memoryInterface_wData :
    io_memoryInterface_memReadData_2; // @[UpdateUnit.scala 68:33]
  wire [127:0] _cacheWriteData_3_T_1 = io_memoryInterface_blockOffset == 2'h3 ? io_memoryInterface_wData :
    io_memoryInterface_memReadData_3; // @[UpdateUnit.scala 68:33]
  wire [127:0] _GEN_1 = io_memoryInterface_rw ? _cacheWriteData_0_T_1 : io_memoryInterface_memReadData_0; // @[UpdateUnit.scala 64:33 68:27 72:22]
  wire [127:0] _GEN_2 = io_memoryInterface_rw ? _cacheWriteData_1_T_1 : io_memoryInterface_memReadData_1; // @[UpdateUnit.scala 64:33 68:27 72:22]
  wire [127:0] _GEN_3 = io_memoryInterface_rw ? _cacheWriteData_2_T_1 : io_memoryInterface_memReadData_2; // @[UpdateUnit.scala 64:33 68:27 72:22]
  wire [127:0] _GEN_4 = io_memoryInterface_rw ? _cacheWriteData_3_T_1 : io_memoryInterface_memReadData_3; // @[UpdateUnit.scala 64:33 68:27 72:22]
  wire [127:0] _GEN_6 = 2'h1 == io_memoryInterface_blockOffset ? io_memoryInterface_memReadData_1 :
    io_memoryInterface_memReadData_0; // @[UpdateUnit.scala 75:{15,15}]
  wire [127:0] _GEN_7 = 2'h2 == io_memoryInterface_blockOffset ? io_memoryInterface_memReadData_2 : _GEN_6; // @[UpdateUnit.scala 75:{15,15}]
  wire [127:0] _GEN_8 = 2'h3 == io_memoryInterface_blockOffset ? io_memoryInterface_memReadData_3 : _GEN_7; // @[UpdateUnit.scala 75:{15,15}]
  wire [127:0] _cacheWriteData_0_T_3 = io_readStage_blockOffset == 2'h0 ? io_readStage_wData :
    io_readStage_memReadData_0; // @[UpdateUnit.scala 89:33]
  wire [127:0] _cacheWriteData_1_T_3 = io_readStage_blockOffset == 2'h1 ? io_readStage_wData :
    io_readStage_memReadData_1; // @[UpdateUnit.scala 89:33]
  wire [127:0] _cacheWriteData_2_T_3 = io_readStage_blockOffset == 2'h2 ? io_readStage_wData :
    io_readStage_memReadData_2; // @[UpdateUnit.scala 89:33]
  wire [127:0] _cacheWriteData_3_T_3 = io_readStage_blockOffset == 2'h3 ? io_readStage_wData :
    io_readStage_memReadData_3; // @[UpdateUnit.scala 89:33]
  wire [127:0] _GEN_10 = io_readStage_rw ? _cacheWriteData_0_T_3 : 128'h0; // @[UpdateUnit.scala 84:27 89:27 53:31]
  wire [127:0] _GEN_11 = io_readStage_rw ? _cacheWriteData_1_T_3 : 128'h0; // @[UpdateUnit.scala 84:27 89:27 53:31]
  wire [127:0] _GEN_12 = io_readStage_rw ? _cacheWriteData_2_T_3 : 128'h0; // @[UpdateUnit.scala 84:27 89:27 53:31]
  wire [127:0] _GEN_13 = io_readStage_rw ? _cacheWriteData_3_T_3 : 128'h0; // @[UpdateUnit.scala 84:27 89:27 53:31]
  wire [127:0] _GEN_15 = 2'h1 == io_readStage_blockOffset ? io_readStage_memReadData_1 : io_readStage_memReadData_0; // @[UpdateUnit.scala 93:{15,15}]
  wire [127:0] _GEN_16 = 2'h2 == io_readStage_blockOffset ? io_readStage_memReadData_2 : _GEN_15; // @[UpdateUnit.scala 93:{15,15}]
  wire [127:0] _GEN_17 = 2'h3 == io_readStage_blockOffset ? io_readStage_memReadData_3 : _GEN_16; // @[UpdateUnit.scala 93:{15,15}]
  wire [3:0] _GEN_18 = io_readStage_valid ? io_readStage_tag : 4'h0; // @[UpdateUnit.scala 42:24 79:34 80:9]
  wire [4:0] _GEN_19 = io_readStage_valid ? io_readStage_index : 5'h0; // @[UpdateUnit.scala 79:34 81:11 43:26]
  wire [2:0] _GEN_20 = io_readStage_valid ? io_readStage_wWay : 3'h0; // @[UpdateUnit.scala 44:24 79:34 82:9]
  wire  _GEN_21 = io_readStage_valid & io_readStage_rw; // @[UpdateUnit.scala 46:27 79:34]
  wire [127:0] _GEN_22 = io_readStage_valid ? _GEN_10 : 128'h0; // @[UpdateUnit.scala 53:31 79:34]
  wire [127:0] _GEN_23 = io_readStage_valid ? _GEN_11 : 128'h0; // @[UpdateUnit.scala 53:31 79:34]
  wire [127:0] _GEN_24 = io_readStage_valid ? _GEN_12 : 128'h0; // @[UpdateUnit.scala 53:31 79:34]
  wire [127:0] _GEN_25 = io_readStage_valid ? _GEN_13 : 128'h0; // @[UpdateUnit.scala 53:31 79:34]
  wire [127:0] _GEN_26 = io_readStage_valid ? _GEN_17 : 128'h0; // @[UpdateUnit.scala 79:34 93:15 50:30]
  wire [1:0] _GEN_27 = io_readStage_valid ? io_readStage_reqId : 2'h0; // @[UpdateUnit.scala 79:34 94:15 49:30]
  wire [1:0] _GEN_28 = io_readStage_valid ? io_readStage_coreId : 2'h0; // @[UpdateUnit.scala 79:34 95:12 48:27]
  wire [4:0] _GEN_32 = io_memoryInterface_valid ? io_memoryInterface_index : _GEN_19; // @[UpdateUnit.scala 57:34 60:11]
  assign io_cacheUpdateControl_tag = io_memoryInterface_valid ? io_memoryInterface_tag : _GEN_18; // @[UpdateUnit.scala 57:34 59:9]
  assign io_cacheUpdateControl_index = _GEN_32[2:0]; // @[UpdateUnit.scala 43:26]
  assign io_cacheUpdateControl_coreId = io_memoryInterface_valid ? io_memoryInterface_coreId : _GEN_28; // @[UpdateUnit.scala 57:34 77:12]
  assign io_cacheUpdateControl_way = io_memoryInterface_valid ? io_memoryInterface_wWay : _GEN_20; // @[UpdateUnit.scala 57:34 61:9]
  assign io_cacheUpdateControl_refill = io_memoryInterface_valid; // @[UpdateUnit.scala 57:34 58:12 45:27]
  assign io_cacheUpdateControl_update = io_memoryInterface_valid ? io_memoryInterface_rw : _GEN_21; // @[UpdateUnit.scala 57:34]
  assign io_cacheUpdateControl_stall = io_memoryInterface_valid & io_readStage_valid; // @[UpdateUnit.scala 99:34]
  assign io_cacheUpdateControl_memWriteData_0 = io_memoryInterface_valid ? _GEN_1 : _GEN_22; // @[UpdateUnit.scala 57:34]
  assign io_cacheUpdateControl_memWriteData_1 = io_memoryInterface_valid ? _GEN_2 : _GEN_23; // @[UpdateUnit.scala 57:34]
  assign io_cacheUpdateControl_memWriteData_2 = io_memoryInterface_valid ? _GEN_3 : _GEN_24; // @[UpdateUnit.scala 57:34]
  assign io_cacheUpdateControl_memWriteData_3 = io_memoryInterface_valid ? _GEN_4 : _GEN_25; // @[UpdateUnit.scala 57:34]
  assign io_cacheUpdateControl_wrEn = io_memoryInterface_valid | _GEN_21; // @[UpdateUnit.scala 57:34 62:10]
  assign io_coreResp_reqId_valid = io_readStage_valid | io_memoryInterface_valid; // @[UpdateUnit.scala 113:49]
  assign io_coreResp_reqId_bits = io_memoryInterface_valid ? io_memoryInterface_reqId : _GEN_27; // @[UpdateUnit.scala 57:34 76:15]
  assign io_coreResp_rData = io_memoryInterface_valid ? _GEN_8 : _GEN_26; // @[UpdateUnit.scala 57:34 75:15]
  assign io_coreResp_responseStatus = io_memoryInterface_valid ? io_memoryInterface_responseStatus : io_readStage_valid; // @[UpdateUnit.scala 57:34 78:20]
endmodule
module RRArbiter(
  input        clock,
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [1:0] io_in_0_bits,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [1:0] io_in_1_bits,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input  [1:0] io_in_2_bits,
  output       io_in_3_ready,
  input        io_in_3_valid,
  input  [1:0] io_in_3_bits,
  input        io_out_ready,
  output       io_out_valid,
  output [1:0] io_out_bits,
  output [1:0] io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 55:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 55:{16,16}]
  wire [1:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits : io_in_0_bits; // @[Arbiter.scala 56:{15,15}]
  wire [1:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits : _GEN_5; // @[Arbiter.scala 56:{15,15}]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [1:0] lastGrant; // @[Reg.scala 19:16]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbiter.scala 81:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbiter.scala 81:49]
  wire  grantMask_3 = 2'h3 > lastGrant; // @[Arbiter.scala 81:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 82:76]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 82:76]
  wire  validMask_3 = io_in_3_valid & grantMask_3; // @[Arbiter.scala 82:76]
  wire  ctrl_2 = ~validMask_1; // @[Arbiter.scala 45:78]
  wire  ctrl_3 = ~(validMask_1 | validMask_2); // @[Arbiter.scala 45:78]
  wire  ctrl_4 = ~(validMask_1 | validMask_2 | validMask_3); // @[Arbiter.scala 45:78]
  wire  ctrl_5 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid); // @[Arbiter.scala 45:78]
  wire  ctrl_6 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 45:78]
  wire  ctrl_7 = ~(validMask_1 | validMask_2 | validMask_3 | io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 45:78]
  wire  _T_3 = grantMask_1 | ctrl_5; // @[Arbiter.scala 86:50]
  wire  _T_5 = ctrl_2 & grantMask_2 | ctrl_6; // @[Arbiter.scala 86:50]
  wire  _T_7 = ctrl_3 & grantMask_3 | ctrl_7; // @[Arbiter.scala 86:50]
  wire [1:0] _GEN_9 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 91:{26,35} 89:41]
  wire [1:0] _GEN_10 = io_in_1_valid ? 2'h1 : _GEN_9; // @[Arbiter.scala 91:{26,35}]
  wire [1:0] _GEN_11 = io_in_0_valid ? 2'h0 : _GEN_10; // @[Arbiter.scala 91:{26,35}]
  wire [1:0] _GEN_12 = validMask_3 ? 2'h3 : _GEN_11; // @[Arbiter.scala 93:{24,33}]
  wire [1:0] _GEN_13 = validMask_2 ? 2'h2 : _GEN_12; // @[Arbiter.scala 93:{24,33}]
  assign io_in_0_ready = ctrl_4 & io_out_ready; // @[Arbiter.scala 74:21]
  assign io_in_1_ready = _T_3 & io_out_ready; // @[Arbiter.scala 74:21]
  assign io_in_2_ready = _T_5 & io_out_ready; // @[Arbiter.scala 74:21]
  assign io_in_3_ready = _T_7 & io_out_ready; // @[Arbiter.scala 74:21]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 55:{16,16}]
  assign io_out_bits = 2'h3 == io_chosen ? io_in_3_bits : _GEN_6; // @[Arbiter.scala 56:{15,15}]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_13; // @[Arbiter.scala 93:{24,33}]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 20:18]
      lastGrant <= io_chosen; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RequestArbiter(
  input          clock,
  output         io_ports_0_reqId_ready,
  input          io_ports_0_reqId_valid,
  input  [1:0]   io_ports_0_reqId_bits,
  input  [14:0]  io_ports_0_addr,
  input          io_ports_0_rw,
  input  [127:0] io_ports_0_wData,
  output         io_ports_1_reqId_ready,
  input          io_ports_1_reqId_valid,
  input  [1:0]   io_ports_1_reqId_bits,
  input  [14:0]  io_ports_1_addr,
  input          io_ports_1_rw,
  input  [127:0] io_ports_1_wData,
  output         io_ports_2_reqId_ready,
  input          io_ports_2_reqId_valid,
  input  [1:0]   io_ports_2_reqId_bits,
  input  [14:0]  io_ports_2_addr,
  input          io_ports_2_rw,
  input  [127:0] io_ports_2_wData,
  output         io_ports_3_reqId_ready,
  input          io_ports_3_reqId_valid,
  input  [1:0]   io_ports_3_reqId_bits,
  input  [14:0]  io_ports_3_addr,
  input          io_ports_3_rw,
  input  [127:0] io_ports_3_wData,
  input          io_out_reqId_ready,
  output         io_out_reqId_valid,
  output [1:0]   io_out_reqId_bits,
  output [14:0]  io_out_addr,
  output         io_out_rw,
  output [127:0] io_out_wData,
  output [1:0]   io_chosen
);
  wire  arbiter_clock; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_0_ready; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_0_valid; // @[RequestArbiter.scala 13:23]
  wire [1:0] arbiter_io_in_0_bits; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_1_ready; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_1_valid; // @[RequestArbiter.scala 13:23]
  wire [1:0] arbiter_io_in_1_bits; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_2_ready; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_2_valid; // @[RequestArbiter.scala 13:23]
  wire [1:0] arbiter_io_in_2_bits; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_3_ready; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_in_3_valid; // @[RequestArbiter.scala 13:23]
  wire [1:0] arbiter_io_in_3_bits; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_out_ready; // @[RequestArbiter.scala 13:23]
  wire  arbiter_io_out_valid; // @[RequestArbiter.scala 13:23]
  wire [1:0] arbiter_io_out_bits; // @[RequestArbiter.scala 13:23]
  wire [1:0] arbiter_io_chosen; // @[RequestArbiter.scala 13:23]
  wire  _GEN_1 = 2'h1 == arbiter_io_chosen ? io_ports_1_rw : io_ports_0_rw; // @[RequestArbiter.scala 22:{13,13}]
  wire  _GEN_2 = 2'h2 == arbiter_io_chosen ? io_ports_2_rw : _GEN_1; // @[RequestArbiter.scala 22:{13,13}]
  wire [127:0] _GEN_5 = 2'h1 == arbiter_io_chosen ? io_ports_1_wData : io_ports_0_wData; // @[RequestArbiter.scala 23:{16,16}]
  wire [127:0] _GEN_6 = 2'h2 == arbiter_io_chosen ? io_ports_2_wData : _GEN_5; // @[RequestArbiter.scala 23:{16,16}]
  wire [14:0] _GEN_9 = 2'h1 == arbiter_io_chosen ? io_ports_1_addr : io_ports_0_addr; // @[RequestArbiter.scala 24:{15,15}]
  wire [14:0] _GEN_10 = 2'h2 == arbiter_io_chosen ? io_ports_2_addr : _GEN_9; // @[RequestArbiter.scala 24:{15,15}]
  RRArbiter arbiter ( // @[RequestArbiter.scala 13:23]
    .clock(arbiter_clock),
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits(arbiter_io_in_0_bits),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits(arbiter_io_in_1_bits),
    .io_in_2_ready(arbiter_io_in_2_ready),
    .io_in_2_valid(arbiter_io_in_2_valid),
    .io_in_2_bits(arbiter_io_in_2_bits),
    .io_in_3_ready(arbiter_io_in_3_ready),
    .io_in_3_valid(arbiter_io_in_3_valid),
    .io_in_3_bits(arbiter_io_in_3_bits),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits(arbiter_io_out_bits),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_ports_0_reqId_ready = arbiter_io_in_0_ready; // @[RequestArbiter.scala 16:27]
  assign io_ports_1_reqId_ready = arbiter_io_in_1_ready; // @[RequestArbiter.scala 16:27]
  assign io_ports_2_reqId_ready = arbiter_io_in_2_ready; // @[RequestArbiter.scala 16:27]
  assign io_ports_3_reqId_ready = arbiter_io_in_3_ready; // @[RequestArbiter.scala 16:27]
  assign io_out_reqId_valid = arbiter_io_out_valid; // @[RequestArbiter.scala 21:16]
  assign io_out_reqId_bits = arbiter_io_out_bits; // @[RequestArbiter.scala 21:16]
  assign io_out_addr = 2'h3 == arbiter_io_chosen ? io_ports_3_addr : _GEN_10; // @[RequestArbiter.scala 24:{15,15}]
  assign io_out_rw = 2'h3 == arbiter_io_chosen ? io_ports_3_rw : _GEN_2; // @[RequestArbiter.scala 22:{13,13}]
  assign io_out_wData = 2'h3 == arbiter_io_chosen ? io_ports_3_wData : _GEN_6; // @[RequestArbiter.scala 23:{16,16}]
  assign io_chosen = arbiter_io_chosen; // @[RequestArbiter.scala 25:13]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_ports_0_reqId_valid; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_0_bits = io_ports_0_reqId_bits; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_1_valid = io_ports_1_reqId_valid; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_1_bits = io_ports_1_reqId_bits; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_2_valid = io_ports_2_reqId_valid; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_2_bits = io_ports_2_reqId_bits; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_3_valid = io_ports_3_reqId_valid; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_in_3_bits = io_ports_3_reqId_bits; // @[RequestArbiter.scala 16:27]
  assign arbiter_io_out_ready = io_out_reqId_ready; // @[RequestArbiter.scala 21:16]
endmodule
module MemBlock(
  input        clock,
  input  [4:0] io_readAddr,
  input  [4:0] io_writeAddr,
  input  [3:0] io_writeData,
  input        io_wrEn,
  output [3:0] io_readData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] mem [0:31]; // @[MemBlock.scala 29:24]
  wire  mem_readData_MPORT_en; // @[MemBlock.scala 29:24]
  wire [4:0] mem_readData_MPORT_addr; // @[MemBlock.scala 29:24]
  wire [3:0] mem_readData_MPORT_data; // @[MemBlock.scala 29:24]
  wire [3:0] mem_MPORT_data; // @[MemBlock.scala 29:24]
  wire [4:0] mem_MPORT_addr; // @[MemBlock.scala 29:24]
  wire  mem_MPORT_mask; // @[MemBlock.scala 29:24]
  wire  mem_MPORT_en; // @[MemBlock.scala 29:24]
  reg [3:0] mem_readData_MPORT_data_pipe_0;
  reg [3:0] writeDataReg; // @[MemBlock.scala 50:29]
  reg  forwardSelReg; // @[MemBlock.scala 51:30]
  wire [3:0] readData = mem_readData_MPORT_data_pipe_0; // @[MemBlock.scala 28:29 48:12]
  assign mem_readData_MPORT_en = 1'h1;
  assign mem_readData_MPORT_addr = io_readAddr;
  assign mem_readData_MPORT_data = mem[mem_readData_MPORT_addr]; // @[MemBlock.scala 29:24]
  assign mem_MPORT_data = io_writeData;
  assign mem_MPORT_addr = io_writeAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEn;
  assign io_readData = forwardSelReg ? writeDataReg : readData; // @[MemBlock.scala 52:21]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[MemBlock.scala 29:24]
    end
    if (1'h1) begin
      mem_readData_MPORT_data_pipe_0 <= mem_readData_MPORT_data;
    end
    writeDataReg <= io_writeData; // @[MemBlock.scala 50:29]
    forwardSelReg <= io_writeAddr == io_readAddr & io_wrEn; // @[MemBlock.scala 51:62]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_readData_MPORT_data_pipe_0 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writeDataReg = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  forwardSelReg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemBlock_8(
  input          clock,
  input  [4:0]   io_readAddr,
  input  [4:0]   io_writeAddr,
  input  [127:0] io_writeData,
  input          io_wrEn,
  output [127:0] io_readData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem [0:31]; // @[MemBlock.scala 29:24]
  wire  mem_readData_MPORT_en; // @[MemBlock.scala 29:24]
  wire [4:0] mem_readData_MPORT_addr; // @[MemBlock.scala 29:24]
  wire [127:0] mem_readData_MPORT_data; // @[MemBlock.scala 29:24]
  wire [127:0] mem_MPORT_data; // @[MemBlock.scala 29:24]
  wire [4:0] mem_MPORT_addr; // @[MemBlock.scala 29:24]
  wire  mem_MPORT_mask; // @[MemBlock.scala 29:24]
  wire  mem_MPORT_en; // @[MemBlock.scala 29:24]
  reg [127:0] mem_readData_MPORT_data_pipe_0;
  reg [127:0] writeDataReg; // @[MemBlock.scala 50:29]
  reg  forwardSelReg; // @[MemBlock.scala 51:30]
  wire [127:0] readData = mem_readData_MPORT_data_pipe_0; // @[MemBlock.scala 28:29 48:12]
  assign mem_readData_MPORT_en = 1'h1;
  assign mem_readData_MPORT_addr = io_readAddr;
  assign mem_readData_MPORT_data = mem[mem_readData_MPORT_addr]; // @[MemBlock.scala 29:24]
  assign mem_MPORT_data = io_writeData;
  assign mem_MPORT_addr = io_writeAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEn;
  assign io_readData = forwardSelReg ? writeDataReg : readData; // @[MemBlock.scala 52:21]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[MemBlock.scala 29:24]
    end
    if (1'h1) begin
      mem_readData_MPORT_data_pipe_0 <= mem_readData_MPORT_data;
    end
    writeDataReg <= io_writeData; // @[MemBlock.scala 50:29]
    forwardSelReg <= io_writeAddr == io_readAddr & io_wrEn; // @[MemBlock.scala 51:62]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {4{`RANDOM}};
  mem_readData_MPORT_data_pipe_0 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  writeDataReg = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  forwardSelReg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheMemory(
  input          clock,
  input  [4:0]   io_rIndex,
  input  [2:0]   io_rWayIdx,
  input  [4:0]   io_wrIndex,
  input  [2:0]   io_wrWayIdx,
  input          io_wrEn,
  input  [127:0] io_wrData_0,
  input  [127:0] io_wrData_1,
  input  [127:0] io_wrData_2,
  input  [127:0] io_wrData_3,
  output [127:0] io_rData_0,
  output [127:0] io_rData_1,
  output [127:0] io_rData_2,
  output [127:0] io_rData_3
);
  wire  MemBlock_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_1_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_1_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_1_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_1_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_1_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_1_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_2_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_2_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_2_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_2_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_2_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_2_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_3_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_3_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_3_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_3_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_3_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_3_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_4_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_4_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_4_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_4_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_4_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_4_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_5_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_5_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_5_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_5_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_5_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_5_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_6_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_6_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_6_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_6_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_6_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_6_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_7_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_7_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_7_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_7_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_7_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_7_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_8_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_8_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_8_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_8_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_8_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_8_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_9_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_9_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_9_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_9_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_9_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_9_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_10_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_10_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_10_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_10_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_10_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_10_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_11_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_11_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_11_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_11_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_11_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_11_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_12_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_12_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_12_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_12_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_12_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_12_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_13_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_13_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_13_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_13_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_13_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_13_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_14_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_14_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_14_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_14_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_14_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_14_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_15_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_15_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_15_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_15_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_15_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_15_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_16_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_16_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_16_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_16_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_16_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_16_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_17_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_17_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_17_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_17_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_17_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_17_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_18_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_18_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_18_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_18_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_18_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_18_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_19_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_19_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_19_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_19_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_19_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_19_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_20_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_20_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_20_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_20_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_20_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_20_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_21_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_21_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_21_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_21_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_21_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_21_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_22_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_22_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_22_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_22_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_22_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_22_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_23_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_23_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_23_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_23_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_23_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_23_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_24_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_24_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_24_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_24_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_24_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_24_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_25_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_25_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_25_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_25_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_25_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_25_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_26_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_26_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_26_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_26_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_26_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_26_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_27_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_27_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_27_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_27_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_27_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_27_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_28_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_28_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_28_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_28_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_28_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_28_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_29_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_29_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_29_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_29_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_29_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_29_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_30_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_30_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_30_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_30_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_30_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_30_io_readData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_31_clock; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_31_io_readAddr; // @[CacheMemory.scala 23:34]
  wire [4:0] MemBlock_31_io_writeAddr; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_31_io_writeData; // @[CacheMemory.scala 23:34]
  wire  MemBlock_31_io_wrEn; // @[CacheMemory.scala 23:34]
  wire [127:0] MemBlock_31_io_readData; // @[CacheMemory.scala 23:34]
  wire [127:0] _GEN_0 = 3'h0 == io_rWayIdx ? MemBlock_io_readData : 128'h0; // @[CacheMemory.scala 26:22 40:37 41:24]
  wire [127:0] _GEN_1 = 3'h0 == io_rWayIdx ? MemBlock_1_io_readData : 128'h0; // @[CacheMemory.scala 26:22 40:37 41:24]
  wire [127:0] _GEN_2 = 3'h0 == io_rWayIdx ? MemBlock_2_io_readData : 128'h0; // @[CacheMemory.scala 26:22 40:37 41:24]
  wire [127:0] _GEN_3 = 3'h0 == io_rWayIdx ? MemBlock_3_io_readData : 128'h0; // @[CacheMemory.scala 26:22 40:37 41:24]
  wire [127:0] _GEN_4 = 3'h1 == io_rWayIdx ? MemBlock_4_io_readData : _GEN_0; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_5 = 3'h1 == io_rWayIdx ? MemBlock_5_io_readData : _GEN_1; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_6 = 3'h1 == io_rWayIdx ? MemBlock_6_io_readData : _GEN_2; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_7 = 3'h1 == io_rWayIdx ? MemBlock_7_io_readData : _GEN_3; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_8 = 3'h2 == io_rWayIdx ? MemBlock_8_io_readData : _GEN_4; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_9 = 3'h2 == io_rWayIdx ? MemBlock_9_io_readData : _GEN_5; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_10 = 3'h2 == io_rWayIdx ? MemBlock_10_io_readData : _GEN_6; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_11 = 3'h2 == io_rWayIdx ? MemBlock_11_io_readData : _GEN_7; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_12 = 3'h3 == io_rWayIdx ? MemBlock_12_io_readData : _GEN_8; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_13 = 3'h3 == io_rWayIdx ? MemBlock_13_io_readData : _GEN_9; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_14 = 3'h3 == io_rWayIdx ? MemBlock_14_io_readData : _GEN_10; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_15 = 3'h3 == io_rWayIdx ? MemBlock_15_io_readData : _GEN_11; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_16 = 3'h4 == io_rWayIdx ? MemBlock_16_io_readData : _GEN_12; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_17 = 3'h4 == io_rWayIdx ? MemBlock_17_io_readData : _GEN_13; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_18 = 3'h4 == io_rWayIdx ? MemBlock_18_io_readData : _GEN_14; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_19 = 3'h4 == io_rWayIdx ? MemBlock_19_io_readData : _GEN_15; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_20 = 3'h5 == io_rWayIdx ? MemBlock_20_io_readData : _GEN_16; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_21 = 3'h5 == io_rWayIdx ? MemBlock_21_io_readData : _GEN_17; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_22 = 3'h5 == io_rWayIdx ? MemBlock_22_io_readData : _GEN_18; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_23 = 3'h5 == io_rWayIdx ? MemBlock_23_io_readData : _GEN_19; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_24 = 3'h6 == io_rWayIdx ? MemBlock_24_io_readData : _GEN_20; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_25 = 3'h6 == io_rWayIdx ? MemBlock_25_io_readData : _GEN_21; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_26 = 3'h6 == io_rWayIdx ? MemBlock_26_io_readData : _GEN_22; // @[CacheMemory.scala 40:37 41:24]
  wire [127:0] _GEN_27 = 3'h6 == io_rWayIdx ? MemBlock_27_io_readData : _GEN_23; // @[CacheMemory.scala 40:37 41:24]
  MemBlock_8 MemBlock ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_clock),
    .io_readAddr(MemBlock_io_readAddr),
    .io_writeAddr(MemBlock_io_writeAddr),
    .io_writeData(MemBlock_io_writeData),
    .io_wrEn(MemBlock_io_wrEn),
    .io_readData(MemBlock_io_readData)
  );
  MemBlock_8 MemBlock_1 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_1_clock),
    .io_readAddr(MemBlock_1_io_readAddr),
    .io_writeAddr(MemBlock_1_io_writeAddr),
    .io_writeData(MemBlock_1_io_writeData),
    .io_wrEn(MemBlock_1_io_wrEn),
    .io_readData(MemBlock_1_io_readData)
  );
  MemBlock_8 MemBlock_2 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_2_clock),
    .io_readAddr(MemBlock_2_io_readAddr),
    .io_writeAddr(MemBlock_2_io_writeAddr),
    .io_writeData(MemBlock_2_io_writeData),
    .io_wrEn(MemBlock_2_io_wrEn),
    .io_readData(MemBlock_2_io_readData)
  );
  MemBlock_8 MemBlock_3 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_3_clock),
    .io_readAddr(MemBlock_3_io_readAddr),
    .io_writeAddr(MemBlock_3_io_writeAddr),
    .io_writeData(MemBlock_3_io_writeData),
    .io_wrEn(MemBlock_3_io_wrEn),
    .io_readData(MemBlock_3_io_readData)
  );
  MemBlock_8 MemBlock_4 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_4_clock),
    .io_readAddr(MemBlock_4_io_readAddr),
    .io_writeAddr(MemBlock_4_io_writeAddr),
    .io_writeData(MemBlock_4_io_writeData),
    .io_wrEn(MemBlock_4_io_wrEn),
    .io_readData(MemBlock_4_io_readData)
  );
  MemBlock_8 MemBlock_5 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_5_clock),
    .io_readAddr(MemBlock_5_io_readAddr),
    .io_writeAddr(MemBlock_5_io_writeAddr),
    .io_writeData(MemBlock_5_io_writeData),
    .io_wrEn(MemBlock_5_io_wrEn),
    .io_readData(MemBlock_5_io_readData)
  );
  MemBlock_8 MemBlock_6 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_6_clock),
    .io_readAddr(MemBlock_6_io_readAddr),
    .io_writeAddr(MemBlock_6_io_writeAddr),
    .io_writeData(MemBlock_6_io_writeData),
    .io_wrEn(MemBlock_6_io_wrEn),
    .io_readData(MemBlock_6_io_readData)
  );
  MemBlock_8 MemBlock_7 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_7_clock),
    .io_readAddr(MemBlock_7_io_readAddr),
    .io_writeAddr(MemBlock_7_io_writeAddr),
    .io_writeData(MemBlock_7_io_writeData),
    .io_wrEn(MemBlock_7_io_wrEn),
    .io_readData(MemBlock_7_io_readData)
  );
  MemBlock_8 MemBlock_8 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_8_clock),
    .io_readAddr(MemBlock_8_io_readAddr),
    .io_writeAddr(MemBlock_8_io_writeAddr),
    .io_writeData(MemBlock_8_io_writeData),
    .io_wrEn(MemBlock_8_io_wrEn),
    .io_readData(MemBlock_8_io_readData)
  );
  MemBlock_8 MemBlock_9 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_9_clock),
    .io_readAddr(MemBlock_9_io_readAddr),
    .io_writeAddr(MemBlock_9_io_writeAddr),
    .io_writeData(MemBlock_9_io_writeData),
    .io_wrEn(MemBlock_9_io_wrEn),
    .io_readData(MemBlock_9_io_readData)
  );
  MemBlock_8 MemBlock_10 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_10_clock),
    .io_readAddr(MemBlock_10_io_readAddr),
    .io_writeAddr(MemBlock_10_io_writeAddr),
    .io_writeData(MemBlock_10_io_writeData),
    .io_wrEn(MemBlock_10_io_wrEn),
    .io_readData(MemBlock_10_io_readData)
  );
  MemBlock_8 MemBlock_11 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_11_clock),
    .io_readAddr(MemBlock_11_io_readAddr),
    .io_writeAddr(MemBlock_11_io_writeAddr),
    .io_writeData(MemBlock_11_io_writeData),
    .io_wrEn(MemBlock_11_io_wrEn),
    .io_readData(MemBlock_11_io_readData)
  );
  MemBlock_8 MemBlock_12 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_12_clock),
    .io_readAddr(MemBlock_12_io_readAddr),
    .io_writeAddr(MemBlock_12_io_writeAddr),
    .io_writeData(MemBlock_12_io_writeData),
    .io_wrEn(MemBlock_12_io_wrEn),
    .io_readData(MemBlock_12_io_readData)
  );
  MemBlock_8 MemBlock_13 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_13_clock),
    .io_readAddr(MemBlock_13_io_readAddr),
    .io_writeAddr(MemBlock_13_io_writeAddr),
    .io_writeData(MemBlock_13_io_writeData),
    .io_wrEn(MemBlock_13_io_wrEn),
    .io_readData(MemBlock_13_io_readData)
  );
  MemBlock_8 MemBlock_14 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_14_clock),
    .io_readAddr(MemBlock_14_io_readAddr),
    .io_writeAddr(MemBlock_14_io_writeAddr),
    .io_writeData(MemBlock_14_io_writeData),
    .io_wrEn(MemBlock_14_io_wrEn),
    .io_readData(MemBlock_14_io_readData)
  );
  MemBlock_8 MemBlock_15 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_15_clock),
    .io_readAddr(MemBlock_15_io_readAddr),
    .io_writeAddr(MemBlock_15_io_writeAddr),
    .io_writeData(MemBlock_15_io_writeData),
    .io_wrEn(MemBlock_15_io_wrEn),
    .io_readData(MemBlock_15_io_readData)
  );
  MemBlock_8 MemBlock_16 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_16_clock),
    .io_readAddr(MemBlock_16_io_readAddr),
    .io_writeAddr(MemBlock_16_io_writeAddr),
    .io_writeData(MemBlock_16_io_writeData),
    .io_wrEn(MemBlock_16_io_wrEn),
    .io_readData(MemBlock_16_io_readData)
  );
  MemBlock_8 MemBlock_17 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_17_clock),
    .io_readAddr(MemBlock_17_io_readAddr),
    .io_writeAddr(MemBlock_17_io_writeAddr),
    .io_writeData(MemBlock_17_io_writeData),
    .io_wrEn(MemBlock_17_io_wrEn),
    .io_readData(MemBlock_17_io_readData)
  );
  MemBlock_8 MemBlock_18 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_18_clock),
    .io_readAddr(MemBlock_18_io_readAddr),
    .io_writeAddr(MemBlock_18_io_writeAddr),
    .io_writeData(MemBlock_18_io_writeData),
    .io_wrEn(MemBlock_18_io_wrEn),
    .io_readData(MemBlock_18_io_readData)
  );
  MemBlock_8 MemBlock_19 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_19_clock),
    .io_readAddr(MemBlock_19_io_readAddr),
    .io_writeAddr(MemBlock_19_io_writeAddr),
    .io_writeData(MemBlock_19_io_writeData),
    .io_wrEn(MemBlock_19_io_wrEn),
    .io_readData(MemBlock_19_io_readData)
  );
  MemBlock_8 MemBlock_20 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_20_clock),
    .io_readAddr(MemBlock_20_io_readAddr),
    .io_writeAddr(MemBlock_20_io_writeAddr),
    .io_writeData(MemBlock_20_io_writeData),
    .io_wrEn(MemBlock_20_io_wrEn),
    .io_readData(MemBlock_20_io_readData)
  );
  MemBlock_8 MemBlock_21 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_21_clock),
    .io_readAddr(MemBlock_21_io_readAddr),
    .io_writeAddr(MemBlock_21_io_writeAddr),
    .io_writeData(MemBlock_21_io_writeData),
    .io_wrEn(MemBlock_21_io_wrEn),
    .io_readData(MemBlock_21_io_readData)
  );
  MemBlock_8 MemBlock_22 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_22_clock),
    .io_readAddr(MemBlock_22_io_readAddr),
    .io_writeAddr(MemBlock_22_io_writeAddr),
    .io_writeData(MemBlock_22_io_writeData),
    .io_wrEn(MemBlock_22_io_wrEn),
    .io_readData(MemBlock_22_io_readData)
  );
  MemBlock_8 MemBlock_23 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_23_clock),
    .io_readAddr(MemBlock_23_io_readAddr),
    .io_writeAddr(MemBlock_23_io_writeAddr),
    .io_writeData(MemBlock_23_io_writeData),
    .io_wrEn(MemBlock_23_io_wrEn),
    .io_readData(MemBlock_23_io_readData)
  );
  MemBlock_8 MemBlock_24 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_24_clock),
    .io_readAddr(MemBlock_24_io_readAddr),
    .io_writeAddr(MemBlock_24_io_writeAddr),
    .io_writeData(MemBlock_24_io_writeData),
    .io_wrEn(MemBlock_24_io_wrEn),
    .io_readData(MemBlock_24_io_readData)
  );
  MemBlock_8 MemBlock_25 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_25_clock),
    .io_readAddr(MemBlock_25_io_readAddr),
    .io_writeAddr(MemBlock_25_io_writeAddr),
    .io_writeData(MemBlock_25_io_writeData),
    .io_wrEn(MemBlock_25_io_wrEn),
    .io_readData(MemBlock_25_io_readData)
  );
  MemBlock_8 MemBlock_26 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_26_clock),
    .io_readAddr(MemBlock_26_io_readAddr),
    .io_writeAddr(MemBlock_26_io_writeAddr),
    .io_writeData(MemBlock_26_io_writeData),
    .io_wrEn(MemBlock_26_io_wrEn),
    .io_readData(MemBlock_26_io_readData)
  );
  MemBlock_8 MemBlock_27 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_27_clock),
    .io_readAddr(MemBlock_27_io_readAddr),
    .io_writeAddr(MemBlock_27_io_writeAddr),
    .io_writeData(MemBlock_27_io_writeData),
    .io_wrEn(MemBlock_27_io_wrEn),
    .io_readData(MemBlock_27_io_readData)
  );
  MemBlock_8 MemBlock_28 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_28_clock),
    .io_readAddr(MemBlock_28_io_readAddr),
    .io_writeAddr(MemBlock_28_io_writeAddr),
    .io_writeData(MemBlock_28_io_writeData),
    .io_wrEn(MemBlock_28_io_wrEn),
    .io_readData(MemBlock_28_io_readData)
  );
  MemBlock_8 MemBlock_29 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_29_clock),
    .io_readAddr(MemBlock_29_io_readAddr),
    .io_writeAddr(MemBlock_29_io_writeAddr),
    .io_writeData(MemBlock_29_io_writeData),
    .io_wrEn(MemBlock_29_io_wrEn),
    .io_readData(MemBlock_29_io_readData)
  );
  MemBlock_8 MemBlock_30 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_30_clock),
    .io_readAddr(MemBlock_30_io_readAddr),
    .io_writeAddr(MemBlock_30_io_writeAddr),
    .io_writeData(MemBlock_30_io_writeData),
    .io_wrEn(MemBlock_30_io_wrEn),
    .io_readData(MemBlock_30_io_readData)
  );
  MemBlock_8 MemBlock_31 ( // @[CacheMemory.scala 23:34]
    .clock(MemBlock_31_clock),
    .io_readAddr(MemBlock_31_io_readAddr),
    .io_writeAddr(MemBlock_31_io_writeAddr),
    .io_writeData(MemBlock_31_io_writeData),
    .io_wrEn(MemBlock_31_io_wrEn),
    .io_readData(MemBlock_31_io_readData)
  );
  assign io_rData_0 = 3'h7 == io_rWayIdx ? MemBlock_28_io_readData : _GEN_24; // @[CacheMemory.scala 40:37 41:24]
  assign io_rData_1 = 3'h7 == io_rWayIdx ? MemBlock_29_io_readData : _GEN_25; // @[CacheMemory.scala 40:37 41:24]
  assign io_rData_2 = 3'h7 == io_rWayIdx ? MemBlock_30_io_readData : _GEN_26; // @[CacheMemory.scala 40:37 41:24]
  assign io_rData_3 = 3'h7 == io_rWayIdx ? MemBlock_31_io_readData : _GEN_27; // @[CacheMemory.scala 40:37 41:24]
  assign MemBlock_clock = clock;
  assign MemBlock_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_io_wrEn = io_wrEn & 3'h0 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_1_clock = clock;
  assign MemBlock_1_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_1_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_1_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_1_io_wrEn = io_wrEn & 3'h0 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_2_clock = clock;
  assign MemBlock_2_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_2_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_2_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_2_io_wrEn = io_wrEn & 3'h0 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_3_clock = clock;
  assign MemBlock_3_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_3_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_3_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_3_io_wrEn = io_wrEn & 3'h0 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_4_clock = clock;
  assign MemBlock_4_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_4_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_4_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_4_io_wrEn = io_wrEn & 3'h1 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_5_clock = clock;
  assign MemBlock_5_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_5_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_5_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_5_io_wrEn = io_wrEn & 3'h1 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_6_clock = clock;
  assign MemBlock_6_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_6_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_6_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_6_io_wrEn = io_wrEn & 3'h1 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_7_clock = clock;
  assign MemBlock_7_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_7_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_7_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_7_io_wrEn = io_wrEn & 3'h1 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_8_clock = clock;
  assign MemBlock_8_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_8_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_8_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_8_io_wrEn = io_wrEn & 3'h2 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_9_clock = clock;
  assign MemBlock_9_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_9_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_9_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_9_io_wrEn = io_wrEn & 3'h2 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_10_clock = clock;
  assign MemBlock_10_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_10_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_10_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_10_io_wrEn = io_wrEn & 3'h2 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_11_clock = clock;
  assign MemBlock_11_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_11_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_11_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_11_io_wrEn = io_wrEn & 3'h2 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_12_clock = clock;
  assign MemBlock_12_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_12_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_12_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_12_io_wrEn = io_wrEn & 3'h3 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_13_clock = clock;
  assign MemBlock_13_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_13_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_13_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_13_io_wrEn = io_wrEn & 3'h3 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_14_clock = clock;
  assign MemBlock_14_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_14_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_14_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_14_io_wrEn = io_wrEn & 3'h3 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_15_clock = clock;
  assign MemBlock_15_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_15_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_15_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_15_io_wrEn = io_wrEn & 3'h3 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_16_clock = clock;
  assign MemBlock_16_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_16_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_16_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_16_io_wrEn = io_wrEn & 3'h4 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_17_clock = clock;
  assign MemBlock_17_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_17_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_17_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_17_io_wrEn = io_wrEn & 3'h4 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_18_clock = clock;
  assign MemBlock_18_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_18_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_18_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_18_io_wrEn = io_wrEn & 3'h4 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_19_clock = clock;
  assign MemBlock_19_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_19_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_19_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_19_io_wrEn = io_wrEn & 3'h4 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_20_clock = clock;
  assign MemBlock_20_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_20_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_20_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_20_io_wrEn = io_wrEn & 3'h5 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_21_clock = clock;
  assign MemBlock_21_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_21_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_21_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_21_io_wrEn = io_wrEn & 3'h5 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_22_clock = clock;
  assign MemBlock_22_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_22_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_22_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_22_io_wrEn = io_wrEn & 3'h5 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_23_clock = clock;
  assign MemBlock_23_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_23_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_23_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_23_io_wrEn = io_wrEn & 3'h5 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_24_clock = clock;
  assign MemBlock_24_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_24_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_24_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_24_io_wrEn = io_wrEn & 3'h6 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_25_clock = clock;
  assign MemBlock_25_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_25_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_25_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_25_io_wrEn = io_wrEn & 3'h6 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_26_clock = clock;
  assign MemBlock_26_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_26_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_26_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_26_io_wrEn = io_wrEn & 3'h6 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_27_clock = clock;
  assign MemBlock_27_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_27_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_27_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_27_io_wrEn = io_wrEn & 3'h6 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_28_clock = clock;
  assign MemBlock_28_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_28_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_28_io_writeData = io_wrData_0; // @[CacheMemory.scala 35:49]
  assign MemBlock_28_io_wrEn = io_wrEn & 3'h7 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_29_clock = clock;
  assign MemBlock_29_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_29_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_29_io_writeData = io_wrData_1; // @[CacheMemory.scala 35:49]
  assign MemBlock_29_io_wrEn = io_wrEn & 3'h7 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_30_clock = clock;
  assign MemBlock_30_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_30_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_30_io_writeData = io_wrData_2; // @[CacheMemory.scala 35:49]
  assign MemBlock_30_io_wrEn = io_wrEn & 3'h7 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
  assign MemBlock_31_clock = clock;
  assign MemBlock_31_io_readAddr = io_rIndex; // @[CacheMemory.scala 34:48]
  assign MemBlock_31_io_writeAddr = io_wrIndex; // @[CacheMemory.scala 36:49]
  assign MemBlock_31_io_writeData = io_wrData_3; // @[CacheMemory.scala 35:49]
  assign MemBlock_31_io_wrEn = io_wrEn & 3'h7 == io_wrWayIdx; // @[CacheMemory.scala 32:30]
endmodule
module RegFifo_8(
  input          clock,
  input          reset,
  input          io_enq_valid,
  input  [511:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [511:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [511:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [511:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [511:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [511:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [511:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [511:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [511:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  always @(posedge clock) begin
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  memReg_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  memReg_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  memReg_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  memReg_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  memReg_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  memReg_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  memReg_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  memReg_7 = _RAND_7[511:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFifo_10(
  input        clock,
  input        reset,
  input        io_enq_valid,
  input  [4:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [4:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] memReg_0; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_1; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_2; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_3; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_4; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_5; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_6; // @[RegFifo.scala 24:19]
  reg [4:0] memReg_7; // @[RegFifo.scala 24:19]
  reg [2:0] readPtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_2 = readPtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _nextVal_T_2; // @[RegFifo.scala 16:22]
  wire [1:0] op = {io_enq_valid,io_deq_ready}; // @[RegFifo.scala 34:25]
  reg  emptyReg; // @[RegFifo.scala 31:25]
  wire  _T_2 = ~emptyReg; // @[RegFifo.scala 40:12]
  wire  _GEN_23 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[RegFifo.scala 37:14 26:29]
  wire  _GEN_26 = 2'h1 == op ? _T_2 : _GEN_23; // @[RegFifo.scala 37:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_26; // @[RegFifo.scala 37:14 26:29]
  reg [2:0] writePtr; // @[RegFifo.scala 15:25]
  wire [2:0] _nextVal_T_5 = writePtr + 3'h1; // @[RegFifo.scala 16:61]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _nextVal_T_5; // @[RegFifo.scala 16:22]
  reg  fullReg; // @[RegFifo.scala 32:24]
  wire  _T_4 = ~fullReg; // @[RegFifo.scala 47:12]
  wire  _GEN_16 = 2'h3 == op & _T_4; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_20 = 2'h2 == op ? _T_4 : _GEN_16; // @[RegFifo.scala 37:14]
  wire  _GEN_27 = 2'h1 == op ? 1'h0 : _GEN_20; // @[RegFifo.scala 37:14 35:28]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_27; // @[RegFifo.scala 37:14 35:28]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[RegFifo.scala 40:23 42:18 31:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[RegFifo.scala 47:22 49:18 31:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[RegFifo.scala 47:22 50:17 32:24]
  wire  _GEN_8 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[RegFifo.scala 58:24 59:19 61:19]
  wire  _GEN_11 = _T_4 ? _GEN_8 : fullReg; // @[RegFifo.scala 55:22 32:24]
  wire  _GEN_12 = fullReg ? 1'h0 : nextRead == nextWrite; // @[RegFifo.scala 67:23 68:20 70:20]
  wire  _GEN_13 = _T_2 ? 1'h0 : _GEN_11; // @[RegFifo.scala 65:23 66:17]
  wire  _GEN_14 = _T_2 ? _GEN_12 : _GEN_6; // @[RegFifo.scala 65:23]
  wire  _GEN_17 = 2'h3 == op ? _GEN_14 : emptyReg; // @[RegFifo.scala 37:14 31:25]
  wire  _GEN_18 = 2'h3 == op ? _GEN_13 : fullReg; // @[RegFifo.scala 37:14 32:24]
  wire  _GEN_21 = 2'h2 == op ? _GEN_6 : _GEN_17; // @[RegFifo.scala 37:14]
  wire  _GEN_25 = 2'h1 == op ? _GEN_3 : _GEN_21; // @[RegFifo.scala 37:14]
  wire  _GEN_29 = 2'h0 == op ? emptyReg : _GEN_25; // @[RegFifo.scala 37:14 31:25]
  wire [4:0] _GEN_49 = 3'h1 == readPtr ? memReg_1 : memReg_0; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_50 = 3'h2 == readPtr ? memReg_2 : _GEN_49; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_51 = 3'h3 == readPtr ? memReg_3 : _GEN_50; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_52 = 3'h4 == readPtr ? memReg_4 : _GEN_51; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_53 = 3'h5 == readPtr ? memReg_5 : _GEN_52; // @[RegFifo.scala 81:{15,15}]
  wire [4:0] _GEN_54 = 3'h6 == readPtr ? memReg_6 : _GEN_53; // @[RegFifo.scala 81:{15,15}]
  wire [3:0] fullNr = fullReg ? 4'h8 : 4'h0; // @[RegFifo.scala 86:19]
  wire [2:0] _number_T_1 = writePtr - readPtr; // @[RegFifo.scala 87:25]
  wire [3:0] _GEN_56 = {{1'd0}, _number_T_1}; // @[RegFifo.scala 87:35]
  wire [3:0] number = _GEN_56 + fullNr; // @[RegFifo.scala 87:35]
  wire  _T_10 = ~reset; // @[RegFifo.scala 88:9]
  wire  _T_21 = readPtr != writePtr; // @[RegFifo.scala 93:16]
  wire  _T_30 = readPtr == writePtr; // @[RegFifo.scala 99:20]
  wire  _T_33 = ~(readPtr == writePtr); // @[RegFifo.scala 99:11]
  wire  _GEN_57 = _T_21 & _T_10; // @[RegFifo.scala 94:11]
  assign io_deq_valid = ~emptyReg; // @[RegFifo.scala 83:19]
  assign io_deq_bits = 3'h7 == readPtr ? memReg_7 : _GEN_54; // @[RegFifo.scala 81:{15,15}]
  always @(posedge clock) begin
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h0 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_0 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h1 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_1 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h2 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_2 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h3 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_3 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h4 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_4 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h5 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_5 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h6 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_6 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (incrWrite) begin // @[RegFifo.scala 77:17]
      if (3'h7 == writePtr) begin // @[RegFifo.scala 78:22]
        memReg_7 <= io_enq_bits; // @[RegFifo.scala 78:22]
      end
    end
    if (reset) begin // @[RegFifo.scala 15:25]
      readPtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrRead) begin // @[RegFifo.scala 17:16]
      if (readPtr == 3'h7) begin // @[RegFifo.scala 16:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_29; // @[RegFifo.scala 31:{25,25}]
    if (reset) begin // @[RegFifo.scala 15:25]
      writePtr <= 3'h0; // @[RegFifo.scala 15:25]
    end else if (incrWrite) begin // @[RegFifo.scala 17:16]
      if (writePtr == 3'h7) begin // @[RegFifo.scala 16:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[RegFifo.scala 32:24]
      fullReg <= 1'h0; // @[RegFifo.scala 32:24]
    end else if (!(2'h0 == op)) begin // @[RegFifo.scala 37:14]
      if (2'h1 == op) begin // @[RegFifo.scala 37:14]
        if (~emptyReg) begin // @[RegFifo.scala 40:23]
          fullReg <= 1'h0; // @[RegFifo.scala 41:17]
        end
      end else if (2'h2 == op) begin // @[RegFifo.scala 37:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_18;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[RegFifo.scala 88:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(number < 4'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:89 assert(number < (depth + 1).U)\n"); // @[RegFifo.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(number < 4'h9) & _T_10) begin
          $fatal; // @[RegFifo.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(emptyReg & fullReg))) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:91 assert(!(emptyReg && fullReg))\n"); // @[RegFifo.scala 91:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(emptyReg & fullReg)) & _T_10) begin
          $fatal; // @[RegFifo.scala 91:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10 & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:94 assert(emptyReg === false.B)\n"); // @[RegFifo.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 94:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & ~_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:95 assert(fullReg === false.B)\n"); // @[RegFifo.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_4 & (_T_21 & _T_10)) begin
          $fatal; // @[RegFifo.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fullReg & _T_10 & ~(readPtr == writePtr)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:99 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 99:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(readPtr == writePtr) & (fullReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 99:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (emptyReg & _T_10 & _T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegFifo.scala:103 assert(readPtr === writePtr)\n"); // @[RegFifo.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_30 & (emptyReg & _T_10)) begin
          $fatal; // @[RegFifo.scala 103:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_4 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_5 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_6 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_7 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  readPtr = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  emptyReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  writePtr = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  fullReg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBackFifo(
  input          clock,
  input          reset,
  input          io_push,
  input          io_pop,
  input  [3:0]   io_pushEntry_tag,
  input  [4:0]   io_pushEntry_index,
  input  [511:0] io_pushEntry_wbData,
  output [3:0]   io_popEntry_tag,
  output [4:0]   io_popEntry_index,
  output [511:0] io_popEntry_wbData,
  output         io_empty
);
  wire  wbDataFifo_clock; // @[WriteBackFifo.scala 22:26]
  wire  wbDataFifo_reset; // @[WriteBackFifo.scala 22:26]
  wire  wbDataFifo_io_enq_valid; // @[WriteBackFifo.scala 22:26]
  wire [511:0] wbDataFifo_io_enq_bits; // @[WriteBackFifo.scala 22:26]
  wire  wbDataFifo_io_deq_ready; // @[WriteBackFifo.scala 22:26]
  wire  wbDataFifo_io_deq_valid; // @[WriteBackFifo.scala 22:26]
  wire [511:0] wbDataFifo_io_deq_bits; // @[WriteBackFifo.scala 22:26]
  wire  tagFifo_clock; // @[WriteBackFifo.scala 23:23]
  wire  tagFifo_reset; // @[WriteBackFifo.scala 23:23]
  wire  tagFifo_io_enq_ready; // @[WriteBackFifo.scala 23:23]
  wire  tagFifo_io_enq_valid; // @[WriteBackFifo.scala 23:23]
  wire [3:0] tagFifo_io_enq_bits; // @[WriteBackFifo.scala 23:23]
  wire  tagFifo_io_deq_ready; // @[WriteBackFifo.scala 23:23]
  wire  tagFifo_io_deq_valid; // @[WriteBackFifo.scala 23:23]
  wire [3:0] tagFifo_io_deq_bits; // @[WriteBackFifo.scala 23:23]
  wire  indexFifo_clock; // @[WriteBackFifo.scala 24:25]
  wire  indexFifo_reset; // @[WriteBackFifo.scala 24:25]
  wire  indexFifo_io_enq_valid; // @[WriteBackFifo.scala 24:25]
  wire [4:0] indexFifo_io_enq_bits; // @[WriteBackFifo.scala 24:25]
  wire  indexFifo_io_deq_ready; // @[WriteBackFifo.scala 24:25]
  wire  indexFifo_io_deq_valid; // @[WriteBackFifo.scala 24:25]
  wire [4:0] indexFifo_io_deq_bits; // @[WriteBackFifo.scala 24:25]
  RegFifo_8 wbDataFifo ( // @[WriteBackFifo.scala 22:26]
    .clock(wbDataFifo_clock),
    .reset(wbDataFifo_reset),
    .io_enq_valid(wbDataFifo_io_enq_valid),
    .io_enq_bits(wbDataFifo_io_enq_bits),
    .io_deq_ready(wbDataFifo_io_deq_ready),
    .io_deq_valid(wbDataFifo_io_deq_valid),
    .io_deq_bits(wbDataFifo_io_deq_bits)
  );
  RegFifo_5 tagFifo ( // @[WriteBackFifo.scala 23:23]
    .clock(tagFifo_clock),
    .reset(tagFifo_reset),
    .io_enq_ready(tagFifo_io_enq_ready),
    .io_enq_valid(tagFifo_io_enq_valid),
    .io_enq_bits(tagFifo_io_enq_bits),
    .io_deq_ready(tagFifo_io_deq_ready),
    .io_deq_valid(tagFifo_io_deq_valid),
    .io_deq_bits(tagFifo_io_deq_bits)
  );
  RegFifo_10 indexFifo ( // @[WriteBackFifo.scala 24:25]
    .clock(indexFifo_clock),
    .reset(indexFifo_reset),
    .io_enq_valid(indexFifo_io_enq_valid),
    .io_enq_bits(indexFifo_io_enq_bits),
    .io_deq_ready(indexFifo_io_deq_ready),
    .io_deq_valid(indexFifo_io_deq_valid),
    .io_deq_bits(indexFifo_io_deq_bits)
  );
  assign io_popEntry_tag = tagFifo_io_deq_bits; // @[WriteBackFifo.scala 40:19]
  assign io_popEntry_index = indexFifo_io_deq_bits; // @[WriteBackFifo.scala 41:21]
  assign io_popEntry_wbData = wbDataFifo_io_deq_bits; // @[WriteBackFifo.scala 42:22]
  assign io_empty = ~wbDataFifo_io_deq_valid | ~tagFifo_io_deq_valid | ~indexFifo_io_deq_valid; // @[WriteBackFifo.scala 28:70]
  assign wbDataFifo_clock = clock;
  assign wbDataFifo_reset = reset;
  assign wbDataFifo_io_enq_valid = io_push; // @[WriteBackFifo.scala 30:27]
  assign wbDataFifo_io_enq_bits = io_pushEntry_wbData; // @[WriteBackFifo.scala 35:26]
  assign wbDataFifo_io_deq_ready = io_pop; // @[WriteBackFifo.scala 37:27]
  assign tagFifo_clock = clock;
  assign tagFifo_reset = reset;
  assign tagFifo_io_enq_valid = io_push; // @[WriteBackFifo.scala 31:24]
  assign tagFifo_io_enq_bits = io_pushEntry_tag; // @[WriteBackFifo.scala 33:23]
  assign tagFifo_io_deq_ready = io_pop; // @[WriteBackFifo.scala 38:24]
  assign indexFifo_clock = clock;
  assign indexFifo_reset = reset;
  assign indexFifo_io_enq_valid = io_push; // @[WriteBackFifo.scala 32:26]
  assign indexFifo_io_enq_bits = io_pushEntry_index; // @[WriteBackFifo.scala 34:25]
  assign indexFifo_io_deq_ready = io_pop; // @[WriteBackFifo.scala 39:26]
endmodule
module MemoryInterface(
  input          clock,
  input          reset,
  input          io_missFifo_popEntry_rw,
  input  [1:0]   io_missFifo_popEntry_reqId,
  input  [1:0]   io_missFifo_popEntry_coreId,
  input  [127:0] io_missFifo_popEntry_wData,
  input  [2:0]   io_missFifo_popEntry_replaceWay,
  input  [3:0]   io_missFifo_popEntry_tag,
  input  [4:0]   io_missFifo_popEntry_index,
  input  [1:0]   io_missFifo_popEntry_blockOffset,
  input          io_missFifo_empty,
  output         io_missFifo_pop,
  input  [3:0]   io_wbFifo_popEntry_tag,
  input  [4:0]   io_wbFifo_popEntry_index,
  input  [511:0] io_wbFifo_popEntry_wbData,
  input          io_wbFifo_empty,
  output         io_wbFifo_pop,
  output         io_updateLogic_valid,
  output [1:0]   io_updateLogic_reqId,
  output [1:0]   io_updateLogic_coreId,
  output         io_updateLogic_rw,
  output [127:0] io_updateLogic_wData,
  output [2:0]   io_updateLogic_wWay,
  output         io_updateLogic_responseStatus,
  output [3:0]   io_updateLogic_tag,
  output [4:0]   io_updateLogic_index,
  output [1:0]   io_updateLogic_blockOffset,
  output [127:0] io_updateLogic_memReadData_0,
  output [127:0] io_updateLogic_memReadData_1,
  output [127:0] io_updateLogic_memReadData_2,
  output [127:0] io_updateLogic_memReadData_3,
  input          io_memController_rChannel_rAddr_ready,
  output         io_memController_rChannel_rAddr_valid,
  output [14:0]  io_memController_rChannel_rAddr_bits,
  output         io_memController_rChannel_rData_ready,
  input          io_memController_rChannel_rData_valid,
  input  [15:0]  io_memController_rChannel_rData_bits,
  input          io_memController_rChannel_rLast,
  input          io_memController_wChannel_wAddr_ready,
  output         io_memController_wChannel_wAddr_valid,
  output [14:0]  io_memController_wChannel_wAddr_bits,
  input          io_memController_wChannel_wData_ready,
  output         io_memController_wChannel_wData_valid,
  output [15:0]  io_memController_wChannel_wData_bits,
  output         io_memController_wChannel_wLast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg; // @[MemoryInterface.scala 45:25]
  reg [15:0] memRwDataReg_0; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_1; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_2; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_3; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_4; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_5; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_6; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_7; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_8; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_9; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_10; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_11; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_12; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_13; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_14; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_15; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_16; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_17; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_18; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_19; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_20; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_21; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_22; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_23; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_24; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_25; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_26; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_27; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_28; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_29; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_30; // @[MemoryInterface.scala 48:29]
  reg [15:0] memRwDataReg_31; // @[MemoryInterface.scala 48:29]
  reg [4:0] burstCounter; // @[MemoryInterface.scala 49:29]
  reg  reqRwReg; // @[MemoryInterface.scala 50:25]
  reg [127:0] reqWDataReg; // @[MemoryInterface.scala 51:28]
  reg [2:0] reqWayReg; // @[MemoryInterface.scala 52:26]
  reg [1:0] reqBlockOffsetReg; // @[MemoryInterface.scala 53:34]
  reg [4:0] reqIndexReg; // @[MemoryInterface.scala 54:28]
  reg [3:0] reqTagReg; // @[MemoryInterface.scala 55:26]
  reg [1:0] reqIdReg; // @[MemoryInterface.scala 56:25]
  reg [1:0] coreIdReg; // @[MemoryInterface.scala 57:26]
  wire [127:0] memRwDataRegAsUint_lo_lo = {memRwDataReg_7,memRwDataReg_6,memRwDataReg_5,memRwDataReg_4,memRwDataReg_3,
    memRwDataReg_2,memRwDataReg_1,memRwDataReg_0}; // @[MemoryInterface.scala 71:41]
  wire [255:0] memRwDataRegAsUint_lo = {memRwDataReg_15,memRwDataReg_14,memRwDataReg_13,memRwDataReg_12,memRwDataReg_11,
    memRwDataReg_10,memRwDataReg_9,memRwDataReg_8,memRwDataRegAsUint_lo_lo}; // @[MemoryInterface.scala 71:41]
  wire [127:0] memRwDataRegAsUint_hi_lo = {memRwDataReg_23,memRwDataReg_22,memRwDataReg_21,memRwDataReg_20,
    memRwDataReg_19,memRwDataReg_18,memRwDataReg_17,memRwDataReg_16}; // @[MemoryInterface.scala 71:41]
  wire [511:0] memRwDataRegAsUint = {memRwDataReg_31,memRwDataReg_30,memRwDataReg_29,memRwDataReg_28,memRwDataReg_27,
    memRwDataReg_26,memRwDataReg_25,memRwDataReg_24,memRwDataRegAsUint_hi_lo,memRwDataRegAsUint_lo}; // @[MemoryInterface.scala 71:41]
  wire  _GEN_0 = ~io_missFifo_empty ? io_missFifo_popEntry_rw : reqRwReg; // @[MemoryInterface.scala 91:38 93:18 50:25]
  wire  _GEN_41 = ~io_wbFifo_empty | _GEN_0; // @[MemoryInterface.scala 77:30 83:18]
  wire [2:0] _GEN_51 = io_memController_wChannel_wAddr_ready ? 3'h4 : stateReg; // @[MemoryInterface.scala 115:51 116:18 45:25]
  wire [4:0] _burstCounter_T_1 = burstCounter + 5'h1; // @[MemoryInterface.scala 123:38]
  wire [15:0] _GEN_52 = 5'h0 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_0; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_53 = 5'h1 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_1; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_54 = 5'h2 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_2; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_55 = 5'h3 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_3; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_56 = 5'h4 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_4; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_57 = 5'h5 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_5; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_58 = 5'h6 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_6; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_59 = 5'h7 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_7; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_60 = 5'h8 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_8; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_61 = 5'h9 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_9; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_62 = 5'ha == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_10; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_63 = 5'hb == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_11; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_64 = 5'hc == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_12; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_65 = 5'hd == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_13; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_66 = 5'he == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_14; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_67 = 5'hf == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_15; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_68 = 5'h10 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_16; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_69 = 5'h11 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_17; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_70 = 5'h12 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_18; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_71 = 5'h13 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_19; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_72 = 5'h14 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_20; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_73 = 5'h15 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_21; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_74 = 5'h16 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_22; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_75 = 5'h17 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_23; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_76 = 5'h18 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_24; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_77 = 5'h19 == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_25; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_78 = 5'h1a == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_26; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_79 = 5'h1b == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_27; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_80 = 5'h1c == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_28; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_81 = 5'h1d == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_29; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_82 = 5'h1e == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_30; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [15:0] _GEN_83 = 5'h1f == burstCounter ? io_memController_rChannel_rData_bits : memRwDataReg_31; // @[MemoryInterface.scala 125:{36,36} 48:29]
  wire [4:0] _GEN_84 = io_memController_rChannel_rLast ? 5'h0 : _burstCounter_T_1; // @[MemoryInterface.scala 123:22 127:47 128:24]
  wire [2:0] _GEN_85 = io_memController_rChannel_rLast ? 3'h5 : stateReg; // @[MemoryInterface.scala 127:47 129:20 45:25]
  wire [4:0] _GEN_86 = io_memController_rChannel_rData_valid ? _GEN_84 : burstCounter; // @[MemoryInterface.scala 122:51 49:29]
  wire [15:0] _GEN_87 = io_memController_rChannel_rData_valid ? _GEN_52 : memRwDataReg_0; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_88 = io_memController_rChannel_rData_valid ? _GEN_53 : memRwDataReg_1; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_89 = io_memController_rChannel_rData_valid ? _GEN_54 : memRwDataReg_2; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_90 = io_memController_rChannel_rData_valid ? _GEN_55 : memRwDataReg_3; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_91 = io_memController_rChannel_rData_valid ? _GEN_56 : memRwDataReg_4; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_92 = io_memController_rChannel_rData_valid ? _GEN_57 : memRwDataReg_5; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_93 = io_memController_rChannel_rData_valid ? _GEN_58 : memRwDataReg_6; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_94 = io_memController_rChannel_rData_valid ? _GEN_59 : memRwDataReg_7; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_95 = io_memController_rChannel_rData_valid ? _GEN_60 : memRwDataReg_8; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_96 = io_memController_rChannel_rData_valid ? _GEN_61 : memRwDataReg_9; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_97 = io_memController_rChannel_rData_valid ? _GEN_62 : memRwDataReg_10; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_98 = io_memController_rChannel_rData_valid ? _GEN_63 : memRwDataReg_11; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_99 = io_memController_rChannel_rData_valid ? _GEN_64 : memRwDataReg_12; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_100 = io_memController_rChannel_rData_valid ? _GEN_65 : memRwDataReg_13; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_101 = io_memController_rChannel_rData_valid ? _GEN_66 : memRwDataReg_14; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_102 = io_memController_rChannel_rData_valid ? _GEN_67 : memRwDataReg_15; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_103 = io_memController_rChannel_rData_valid ? _GEN_68 : memRwDataReg_16; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_104 = io_memController_rChannel_rData_valid ? _GEN_69 : memRwDataReg_17; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_105 = io_memController_rChannel_rData_valid ? _GEN_70 : memRwDataReg_18; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_106 = io_memController_rChannel_rData_valid ? _GEN_71 : memRwDataReg_19; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_107 = io_memController_rChannel_rData_valid ? _GEN_72 : memRwDataReg_20; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_108 = io_memController_rChannel_rData_valid ? _GEN_73 : memRwDataReg_21; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_109 = io_memController_rChannel_rData_valid ? _GEN_74 : memRwDataReg_22; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_110 = io_memController_rChannel_rData_valid ? _GEN_75 : memRwDataReg_23; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_111 = io_memController_rChannel_rData_valid ? _GEN_76 : memRwDataReg_24; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_112 = io_memController_rChannel_rData_valid ? _GEN_77 : memRwDataReg_25; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_113 = io_memController_rChannel_rData_valid ? _GEN_78 : memRwDataReg_26; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_114 = io_memController_rChannel_rData_valid ? _GEN_79 : memRwDataReg_27; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_115 = io_memController_rChannel_rData_valid ? _GEN_80 : memRwDataReg_28; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_116 = io_memController_rChannel_rData_valid ? _GEN_81 : memRwDataReg_29; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_117 = io_memController_rChannel_rData_valid ? _GEN_82 : memRwDataReg_30; // @[MemoryInterface.scala 122:51 48:29]
  wire [15:0] _GEN_118 = io_memController_rChannel_rData_valid ? _GEN_83 : memRwDataReg_31; // @[MemoryInterface.scala 122:51 48:29]
  wire [2:0] _GEN_119 = io_memController_rChannel_rData_valid ? _GEN_85 : stateReg; // @[MemoryInterface.scala 122:51 45:25]
  wire [15:0] _GEN_121 = 5'h1 == burstCounter ? memRwDataReg_1 : memRwDataReg_0; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_122 = 5'h2 == burstCounter ? memRwDataReg_2 : _GEN_121; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_123 = 5'h3 == burstCounter ? memRwDataReg_3 : _GEN_122; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_124 = 5'h4 == burstCounter ? memRwDataReg_4 : _GEN_123; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_125 = 5'h5 == burstCounter ? memRwDataReg_5 : _GEN_124; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_126 = 5'h6 == burstCounter ? memRwDataReg_6 : _GEN_125; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_127 = 5'h7 == burstCounter ? memRwDataReg_7 : _GEN_126; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_128 = 5'h8 == burstCounter ? memRwDataReg_8 : _GEN_127; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_129 = 5'h9 == burstCounter ? memRwDataReg_9 : _GEN_128; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_130 = 5'ha == burstCounter ? memRwDataReg_10 : _GEN_129; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_131 = 5'hb == burstCounter ? memRwDataReg_11 : _GEN_130; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_132 = 5'hc == burstCounter ? memRwDataReg_12 : _GEN_131; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_133 = 5'hd == burstCounter ? memRwDataReg_13 : _GEN_132; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_134 = 5'he == burstCounter ? memRwDataReg_14 : _GEN_133; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_135 = 5'hf == burstCounter ? memRwDataReg_15 : _GEN_134; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_136 = 5'h10 == burstCounter ? memRwDataReg_16 : _GEN_135; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_137 = 5'h11 == burstCounter ? memRwDataReg_17 : _GEN_136; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_138 = 5'h12 == burstCounter ? memRwDataReg_18 : _GEN_137; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_139 = 5'h13 == burstCounter ? memRwDataReg_19 : _GEN_138; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_140 = 5'h14 == burstCounter ? memRwDataReg_20 : _GEN_139; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_141 = 5'h15 == burstCounter ? memRwDataReg_21 : _GEN_140; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_142 = 5'h16 == burstCounter ? memRwDataReg_22 : _GEN_141; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_143 = 5'h17 == burstCounter ? memRwDataReg_23 : _GEN_142; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_144 = 5'h18 == burstCounter ? memRwDataReg_24 : _GEN_143; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_145 = 5'h19 == burstCounter ? memRwDataReg_25 : _GEN_144; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_146 = 5'h1a == burstCounter ? memRwDataReg_26 : _GEN_145; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_147 = 5'h1b == burstCounter ? memRwDataReg_27 : _GEN_146; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_148 = 5'h1c == burstCounter ? memRwDataReg_28 : _GEN_147; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_149 = 5'h1d == burstCounter ? memRwDataReg_29 : _GEN_148; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_150 = 5'h1e == burstCounter ? memRwDataReg_30 : _GEN_149; // @[MemoryInterface.scala 136:{16,16}]
  wire [15:0] _GEN_151 = 5'h1f == burstCounter ? memRwDataReg_31 : _GEN_150; // @[MemoryInterface.scala 136:{16,16}]
  wire  _T_7 = burstCounter == 5'h1f; // @[MemoryInterface.scala 141:27]
  wire [4:0] _GEN_153 = burstCounter == 5'h1f ? 5'h0 : _burstCounter_T_1; // @[MemoryInterface.scala 139:22 141:48 143:24]
  wire [2:0] _GEN_154 = burstCounter == 5'h1f ? 3'h6 : stateReg; // @[MemoryInterface.scala 141:48 144:20 45:25]
  wire [4:0] _GEN_155 = io_memController_wChannel_wData_ready ? _GEN_153 : burstCounter; // @[MemoryInterface.scala 138:51 49:29]
  wire  _GEN_156 = io_memController_wChannel_wData_ready & _T_7; // @[MemoryInterface.scala 138:51 65:29]
  wire [2:0] _GEN_157 = io_memController_wChannel_wData_ready ? _GEN_154 : stateReg; // @[MemoryInterface.scala 138:51 45:25]
  wire [2:0] _GEN_159 = 3'h6 == stateReg ? 3'h0 : stateReg; // @[MemoryInterface.scala 158:16 74:20 45:25]
  wire [2:0] _GEN_161 = 3'h5 == stateReg ? 3'h0 : _GEN_159; // @[MemoryInterface.scala 153:16 74:20]
  wire  _GEN_162 = 3'h5 == stateReg ? 1'h0 : 3'h6 == stateReg; // @[MemoryInterface.scala 74:20 66:30]
  wire [15:0] _GEN_164 = 3'h4 == stateReg ? _GEN_151 : 16'h0; // @[MemoryInterface.scala 136:16 74:20 64:29]
  wire [4:0] _GEN_165 = 3'h4 == stateReg ? _GEN_155 : burstCounter; // @[MemoryInterface.scala 74:20 49:29]
  wire [2:0] _GEN_167 = 3'h4 == stateReg ? _GEN_157 : _GEN_161; // @[MemoryInterface.scala 74:20]
  wire  _GEN_168 = 3'h4 == stateReg ? 1'h0 : 3'h5 == stateReg; // @[MemoryInterface.scala 74:20 67:32]
  wire  _GEN_169 = 3'h4 == stateReg ? 1'h0 : _GEN_162; // @[MemoryInterface.scala 74:20 66:30]
  wire [4:0] _GEN_171 = 3'h3 == stateReg ? _GEN_86 : _GEN_165; // @[MemoryInterface.scala 74:20]
  wire [15:0] _GEN_172 = 3'h3 == stateReg ? _GEN_87 : memRwDataReg_0; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_173 = 3'h3 == stateReg ? _GEN_88 : memRwDataReg_1; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_174 = 3'h3 == stateReg ? _GEN_89 : memRwDataReg_2; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_175 = 3'h3 == stateReg ? _GEN_90 : memRwDataReg_3; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_176 = 3'h3 == stateReg ? _GEN_91 : memRwDataReg_4; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_177 = 3'h3 == stateReg ? _GEN_92 : memRwDataReg_5; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_178 = 3'h3 == stateReg ? _GEN_93 : memRwDataReg_6; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_179 = 3'h3 == stateReg ? _GEN_94 : memRwDataReg_7; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_180 = 3'h3 == stateReg ? _GEN_95 : memRwDataReg_8; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_181 = 3'h3 == stateReg ? _GEN_96 : memRwDataReg_9; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_182 = 3'h3 == stateReg ? _GEN_97 : memRwDataReg_10; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_183 = 3'h3 == stateReg ? _GEN_98 : memRwDataReg_11; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_184 = 3'h3 == stateReg ? _GEN_99 : memRwDataReg_12; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_185 = 3'h3 == stateReg ? _GEN_100 : memRwDataReg_13; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_186 = 3'h3 == stateReg ? _GEN_101 : memRwDataReg_14; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_187 = 3'h3 == stateReg ? _GEN_102 : memRwDataReg_15; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_188 = 3'h3 == stateReg ? _GEN_103 : memRwDataReg_16; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_189 = 3'h3 == stateReg ? _GEN_104 : memRwDataReg_17; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_190 = 3'h3 == stateReg ? _GEN_105 : memRwDataReg_18; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_191 = 3'h3 == stateReg ? _GEN_106 : memRwDataReg_19; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_192 = 3'h3 == stateReg ? _GEN_107 : memRwDataReg_20; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_193 = 3'h3 == stateReg ? _GEN_108 : memRwDataReg_21; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_194 = 3'h3 == stateReg ? _GEN_109 : memRwDataReg_22; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_195 = 3'h3 == stateReg ? _GEN_110 : memRwDataReg_23; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_196 = 3'h3 == stateReg ? _GEN_111 : memRwDataReg_24; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_197 = 3'h3 == stateReg ? _GEN_112 : memRwDataReg_25; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_198 = 3'h3 == stateReg ? _GEN_113 : memRwDataReg_26; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_199 = 3'h3 == stateReg ? _GEN_114 : memRwDataReg_27; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_200 = 3'h3 == stateReg ? _GEN_115 : memRwDataReg_28; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_201 = 3'h3 == stateReg ? _GEN_116 : memRwDataReg_29; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_202 = 3'h3 == stateReg ? _GEN_117 : memRwDataReg_30; // @[MemoryInterface.scala 74:20 48:29]
  wire [15:0] _GEN_203 = 3'h3 == stateReg ? _GEN_118 : memRwDataReg_31; // @[MemoryInterface.scala 74:20 48:29]
  wire [2:0] _GEN_204 = 3'h3 == stateReg ? _GEN_119 : _GEN_167; // @[MemoryInterface.scala 74:20]
  wire  _GEN_205 = 3'h3 == stateReg ? 1'h0 : 3'h4 == stateReg; // @[MemoryInterface.scala 74:20 63:34]
  wire [15:0] _GEN_206 = 3'h3 == stateReg ? 16'h0 : _GEN_164; // @[MemoryInterface.scala 74:20 64:29]
  wire  _GEN_207 = 3'h3 == stateReg ? 1'h0 : 3'h4 == stateReg & _GEN_156; // @[MemoryInterface.scala 74:20 65:29]
  wire  _GEN_208 = 3'h3 == stateReg ? 1'h0 : _GEN_168; // @[MemoryInterface.scala 74:20 67:32]
  wire  _GEN_209 = 3'h3 == stateReg ? 1'h0 : _GEN_169; // @[MemoryInterface.scala 74:20 66:30]
  wire  _GEN_212 = 3'h2 == stateReg ? 1'h0 : 3'h3 == stateReg; // @[MemoryInterface.scala 74:20 61:34]
  wire  _GEN_246 = 3'h2 == stateReg ? 1'h0 : _GEN_205; // @[MemoryInterface.scala 74:20 63:34]
  wire [15:0] _GEN_247 = 3'h2 == stateReg ? 16'h0 : _GEN_206; // @[MemoryInterface.scala 74:20 64:29]
  wire  _GEN_248 = 3'h2 == stateReg ? 1'h0 : _GEN_207; // @[MemoryInterface.scala 74:20 65:29]
  wire  _GEN_249 = 3'h2 == stateReg ? 1'h0 : _GEN_208; // @[MemoryInterface.scala 74:20 67:32]
  wire  _GEN_250 = 3'h2 == stateReg ? 1'h0 : _GEN_209; // @[MemoryInterface.scala 74:20 66:30]
  wire  _GEN_253 = 3'h1 == stateReg ? 1'h0 : 3'h2 == stateReg; // @[MemoryInterface.scala 74:20 62:34]
  wire  _GEN_254 = 3'h1 == stateReg ? 1'h0 : _GEN_212; // @[MemoryInterface.scala 74:20 61:34]
  wire  _GEN_288 = 3'h1 == stateReg ? 1'h0 : _GEN_246; // @[MemoryInterface.scala 74:20 63:34]
  wire [15:0] _GEN_289 = 3'h1 == stateReg ? 16'h0 : _GEN_247; // @[MemoryInterface.scala 74:20 64:29]
  wire  _GEN_290 = 3'h1 == stateReg ? 1'h0 : _GEN_248; // @[MemoryInterface.scala 74:20 65:29]
  wire  _GEN_291 = 3'h1 == stateReg ? 1'h0 : _GEN_249; // @[MemoryInterface.scala 74:20 67:32]
  wire  _GEN_292 = 3'h1 == stateReg ? 1'h0 : _GEN_250; // @[MemoryInterface.scala 74:20 66:30]
  wire [8:0] _outAddr_T = {reqTagReg,reqIndexReg}; // @[Cat.scala 33:92]
  wire [14:0] _GEN_343 = {_outAddr_T, 6'h0}; // @[MemoryInterface.scala 176:45]
  wire [15:0] outAddr = {{1'd0}, _GEN_343}; // @[MemoryInterface.scala 176:45]
  assign io_missFifo_pop = 3'h0 == stateReg ? 1'h0 : _GEN_291; // @[MemoryInterface.scala 74:20 67:32]
  assign io_wbFifo_pop = 3'h0 == stateReg ? 1'h0 : _GEN_292; // @[MemoryInterface.scala 74:20 66:30]
  assign io_updateLogic_valid = 3'h0 == stateReg ? 1'h0 : _GEN_291; // @[MemoryInterface.scala 74:20 67:32]
  assign io_updateLogic_reqId = reqIdReg; // @[MemoryInterface.scala 173:24]
  assign io_updateLogic_coreId = coreIdReg; // @[MemoryInterface.scala 174:25]
  assign io_updateLogic_rw = reqRwReg; // @[MemoryInterface.scala 166:21]
  assign io_updateLogic_wData = reqWDataReg; // @[MemoryInterface.scala 167:24]
  assign io_updateLogic_wWay = reqWayReg; // @[MemoryInterface.scala 168:23]
  assign io_updateLogic_responseStatus = 3'h0 == stateReg ? 1'h0 : _GEN_291; // @[MemoryInterface.scala 74:20 67:32]
  assign io_updateLogic_tag = reqTagReg; // @[MemoryInterface.scala 172:22]
  assign io_updateLogic_index = reqIndexReg; // @[MemoryInterface.scala 171:24]
  assign io_updateLogic_blockOffset = reqBlockOffsetReg; // @[MemoryInterface.scala 170:30]
  assign io_updateLogic_memReadData_0 = memRwDataRegAsUint[127:0]; // @[MemoryInterface.scala 179:56]
  assign io_updateLogic_memReadData_1 = memRwDataRegAsUint[255:128]; // @[MemoryInterface.scala 179:56]
  assign io_updateLogic_memReadData_2 = memRwDataRegAsUint[383:256]; // @[MemoryInterface.scala 179:56]
  assign io_updateLogic_memReadData_3 = memRwDataRegAsUint[511:384]; // @[MemoryInterface.scala 179:56]
  assign io_memController_rChannel_rAddr_valid = 3'h0 == stateReg ? 1'h0 : 3'h1 == stateReg; // @[MemoryInterface.scala 74:20 60:34]
  assign io_memController_rChannel_rAddr_bits = outAddr[14:0]; // @[MemoryInterface.scala 183:40]
  assign io_memController_rChannel_rData_ready = 3'h0 == stateReg ? 1'h0 : _GEN_254; // @[MemoryInterface.scala 74:20 61:34]
  assign io_memController_wChannel_wAddr_valid = 3'h0 == stateReg ? 1'h0 : _GEN_253; // @[MemoryInterface.scala 74:20 62:34]
  assign io_memController_wChannel_wAddr_bits = outAddr[14:0]; // @[MemoryInterface.scala 186:40]
  assign io_memController_wChannel_wData_valid = 3'h0 == stateReg ? 1'h0 : _GEN_288; // @[MemoryInterface.scala 74:20 63:34]
  assign io_memController_wChannel_wData_bits = 3'h0 == stateReg ? 16'h0 : _GEN_289; // @[MemoryInterface.scala 74:20 64:29]
  assign io_memController_wChannel_wLast = 3'h0 == stateReg ? 1'h0 : _GEN_290; // @[MemoryInterface.scala 74:20 65:29]
  always @(posedge clock) begin
    if (reset) begin // @[MemoryInterface.scala 45:25]
      stateReg <= 3'h0; // @[MemoryInterface.scala 45:25]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        stateReg <= 3'h2; // @[MemoryInterface.scala 90:18]
      end else if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
        stateReg <= 3'h1; // @[MemoryInterface.scala 102:18]
      end
    end else if (3'h1 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (io_memController_rChannel_rAddr_ready) begin // @[MemoryInterface.scala 108:51]
        stateReg <= 3'h3; // @[MemoryInterface.scala 109:18]
      end
    end else if (3'h2 == stateReg) begin // @[MemoryInterface.scala 74:20]
      stateReg <= _GEN_51;
    end else begin
      stateReg <= _GEN_204;
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_0 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_0 <= io_wbFifo_popEntry_wbData[15:0]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_0 <= _GEN_172;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_1 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_1 <= io_wbFifo_popEntry_wbData[31:16]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_1 <= _GEN_173;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_2 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_2 <= io_wbFifo_popEntry_wbData[47:32]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_2 <= _GEN_174;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_3 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_3 <= io_wbFifo_popEntry_wbData[63:48]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_3 <= _GEN_175;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_4 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_4 <= io_wbFifo_popEntry_wbData[79:64]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_4 <= _GEN_176;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_5 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_5 <= io_wbFifo_popEntry_wbData[95:80]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_5 <= _GEN_177;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_6 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_6 <= io_wbFifo_popEntry_wbData[111:96]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_6 <= _GEN_178;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_7 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_7 <= io_wbFifo_popEntry_wbData[127:112]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_7 <= _GEN_179;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_8 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_8 <= io_wbFifo_popEntry_wbData[143:128]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_8 <= _GEN_180;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_9 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_9 <= io_wbFifo_popEntry_wbData[159:144]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_9 <= _GEN_181;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_10 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_10 <= io_wbFifo_popEntry_wbData[175:160]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_10 <= _GEN_182;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_11 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_11 <= io_wbFifo_popEntry_wbData[191:176]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_11 <= _GEN_183;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_12 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_12 <= io_wbFifo_popEntry_wbData[207:192]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_12 <= _GEN_184;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_13 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_13 <= io_wbFifo_popEntry_wbData[223:208]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_13 <= _GEN_185;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_14 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_14 <= io_wbFifo_popEntry_wbData[239:224]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_14 <= _GEN_186;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_15 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_15 <= io_wbFifo_popEntry_wbData[255:240]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_15 <= _GEN_187;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_16 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_16 <= io_wbFifo_popEntry_wbData[271:256]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_16 <= _GEN_188;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_17 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_17 <= io_wbFifo_popEntry_wbData[287:272]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_17 <= _GEN_189;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_18 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_18 <= io_wbFifo_popEntry_wbData[303:288]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_18 <= _GEN_190;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_19 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_19 <= io_wbFifo_popEntry_wbData[319:304]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_19 <= _GEN_191;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_20 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_20 <= io_wbFifo_popEntry_wbData[335:320]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_20 <= _GEN_192;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_21 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_21 <= io_wbFifo_popEntry_wbData[351:336]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_21 <= _GEN_193;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_22 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_22 <= io_wbFifo_popEntry_wbData[367:352]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_22 <= _GEN_194;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_23 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_23 <= io_wbFifo_popEntry_wbData[383:368]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_23 <= _GEN_195;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_24 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_24 <= io_wbFifo_popEntry_wbData[399:384]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_24 <= _GEN_196;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_25 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_25 <= io_wbFifo_popEntry_wbData[415:400]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_25 <= _GEN_197;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_26 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_26 <= io_wbFifo_popEntry_wbData[431:416]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_26 <= _GEN_198;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_27 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_27 <= io_wbFifo_popEntry_wbData[447:432]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_27 <= _GEN_199;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_28 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_28 <= io_wbFifo_popEntry_wbData[463:448]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_28 <= _GEN_200;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_29 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_29 <= io_wbFifo_popEntry_wbData[479:464]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_29 <= _GEN_201;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_30 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_30 <= io_wbFifo_popEntry_wbData[495:480]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_30 <= _GEN_202;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 48:29]
      memRwDataReg_31 <= 16'h0; // @[MemoryInterface.scala 48:29]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        memRwDataReg_31 <= io_wbFifo_popEntry_wbData[511:496]; // @[MemoryInterface.scala 80:27]
      end
    end else if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        memRwDataReg_31 <= _GEN_203;
      end
    end
    if (reset) begin // @[MemoryInterface.scala 49:29]
      burstCounter <= 5'h0; // @[MemoryInterface.scala 49:29]
    end else if (!(3'h0 == stateReg)) begin // @[MemoryInterface.scala 74:20]
      if (!(3'h1 == stateReg)) begin // @[MemoryInterface.scala 74:20]
        if (!(3'h2 == stateReg)) begin // @[MemoryInterface.scala 74:20]
          burstCounter <= _GEN_171;
        end
      end
    end
    if (reset) begin // @[MemoryInterface.scala 50:25]
      reqRwReg <= 1'h0; // @[MemoryInterface.scala 50:25]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      reqRwReg <= _GEN_41;
    end
    if (reset) begin // @[MemoryInterface.scala 51:28]
      reqWDataReg <= 128'h0; // @[MemoryInterface.scala 51:28]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        reqWDataReg <= 128'h0; // @[MemoryInterface.scala 84:21]
      end else if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
        reqWDataReg <= io_missFifo_popEntry_wData; // @[MemoryInterface.scala 94:21]
      end
    end
    if (reset) begin // @[MemoryInterface.scala 52:26]
      reqWayReg <= 3'h0; // @[MemoryInterface.scala 52:26]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        reqWayReg <= 3'h0; // @[MemoryInterface.scala 85:19]
      end else if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
        reqWayReg <= io_missFifo_popEntry_replaceWay; // @[MemoryInterface.scala 95:19]
      end
    end
    if (reset) begin // @[MemoryInterface.scala 53:34]
      reqBlockOffsetReg <= 2'h0; // @[MemoryInterface.scala 53:34]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        reqBlockOffsetReg <= 2'h0; // @[MemoryInterface.scala 86:27]
      end else if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
        reqBlockOffsetReg <= io_missFifo_popEntry_blockOffset; // @[MemoryInterface.scala 96:27]
      end
    end
    if (reset) begin // @[MemoryInterface.scala 54:28]
      reqIndexReg <= 5'h0; // @[MemoryInterface.scala 54:28]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        reqIndexReg <= io_wbFifo_popEntry_index; // @[MemoryInterface.scala 87:21]
      end else if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
        reqIndexReg <= io_missFifo_popEntry_index; // @[MemoryInterface.scala 97:21]
      end
    end
    if (reset) begin // @[MemoryInterface.scala 55:26]
      reqTagReg <= 4'h0; // @[MemoryInterface.scala 55:26]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (~io_wbFifo_empty) begin // @[MemoryInterface.scala 77:30]
        reqTagReg <= io_wbFifo_popEntry_tag; // @[MemoryInterface.scala 88:19]
      end else if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
        reqTagReg <= io_missFifo_popEntry_tag; // @[MemoryInterface.scala 98:19]
      end
    end
    if (reset) begin // @[MemoryInterface.scala 56:25]
      reqIdReg <= 2'h0; // @[MemoryInterface.scala 56:25]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (!(~io_wbFifo_empty)) begin // @[MemoryInterface.scala 77:30]
        if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
          reqIdReg <= io_missFifo_popEntry_reqId; // @[MemoryInterface.scala 99:18]
        end
      end
    end
    if (reset) begin // @[MemoryInterface.scala 57:26]
      coreIdReg <= 2'h0; // @[MemoryInterface.scala 57:26]
    end else if (3'h0 == stateReg) begin // @[MemoryInterface.scala 74:20]
      if (!(~io_wbFifo_empty)) begin // @[MemoryInterface.scala 77:30]
        if (~io_missFifo_empty) begin // @[MemoryInterface.scala 91:38]
          coreIdReg <= io_missFifo_popEntry_coreId; // @[MemoryInterface.scala 100:19]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  memRwDataReg_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  memRwDataReg_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  memRwDataReg_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  memRwDataReg_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  memRwDataReg_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  memRwDataReg_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  memRwDataReg_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  memRwDataReg_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  memRwDataReg_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  memRwDataReg_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  memRwDataReg_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  memRwDataReg_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  memRwDataReg_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  memRwDataReg_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  memRwDataReg_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  memRwDataReg_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  memRwDataReg_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  memRwDataReg_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  memRwDataReg_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  memRwDataReg_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  memRwDataReg_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  memRwDataReg_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  memRwDataReg_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  memRwDataReg_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  memRwDataReg_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  memRwDataReg_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  memRwDataReg_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  memRwDataReg_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  memRwDataReg_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  memRwDataReg_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  memRwDataReg_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  memRwDataReg_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  burstCounter = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  reqRwReg = _RAND_34[0:0];
  _RAND_35 = {4{`RANDOM}};
  reqWDataReg = _RAND_35[127:0];
  _RAND_36 = {1{`RANDOM}};
  reqWayReg = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  reqBlockOffsetReg = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  reqIndexReg = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  reqTagReg = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  reqIdReg = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  coreIdReg = _RAND_41[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SharedPipelinedCache(
  input          clock,
  input          reset,
  output         io_cache_coreReqs_0_reqId_ready,
  input          io_cache_coreReqs_0_reqId_valid,
  input  [1:0]   io_cache_coreReqs_0_reqId_bits,
  input  [14:0]  io_cache_coreReqs_0_addr,
  input          io_cache_coreReqs_0_rw,
  input  [127:0] io_cache_coreReqs_0_wData,
  output         io_cache_coreReqs_1_reqId_ready,
  input          io_cache_coreReqs_1_reqId_valid,
  input  [1:0]   io_cache_coreReqs_1_reqId_bits,
  input  [14:0]  io_cache_coreReqs_1_addr,
  input          io_cache_coreReqs_1_rw,
  input  [127:0] io_cache_coreReqs_1_wData,
  output         io_cache_coreReqs_2_reqId_ready,
  input          io_cache_coreReqs_2_reqId_valid,
  input  [1:0]   io_cache_coreReqs_2_reqId_bits,
  input  [14:0]  io_cache_coreReqs_2_addr,
  input          io_cache_coreReqs_2_rw,
  input  [127:0] io_cache_coreReqs_2_wData,
  output         io_cache_coreReqs_3_reqId_ready,
  input          io_cache_coreReqs_3_reqId_valid,
  input  [1:0]   io_cache_coreReqs_3_reqId_bits,
  input  [14:0]  io_cache_coreReqs_3_addr,
  input          io_cache_coreReqs_3_rw,
  input  [127:0] io_cache_coreReqs_3_wData,
  output         io_cache_coreResps_0_reqId_valid,
  output [1:0]   io_cache_coreResps_0_reqId_bits,
  output [127:0] io_cache_coreResps_0_rData,
  output         io_cache_coreResps_0_responseStatus,
  output         io_cache_coreResps_1_reqId_valid,
  output [1:0]   io_cache_coreResps_1_reqId_bits,
  output [127:0] io_cache_coreResps_1_rData,
  output         io_cache_coreResps_1_responseStatus,
  output         io_cache_coreResps_2_reqId_valid,
  output [1:0]   io_cache_coreResps_2_reqId_bits,
  output [127:0] io_cache_coreResps_2_rData,
  output         io_cache_coreResps_2_responseStatus,
  output         io_cache_coreResps_3_reqId_valid,
  output [1:0]   io_cache_coreResps_3_reqId_bits,
  output [127:0] io_cache_coreResps_3_rData,
  output         io_cache_coreResps_3_responseStatus,
  output         io_repPol_update_valid,
  output [2:0]   io_repPol_update_bits,
  output         io_repPol_stall,
  output [4:0]   io_repPol_setIdx,
  input  [2:0]   io_repPol_replaceWay,
  input          io_mem_rChannel_rAddr_ready,
  output         io_mem_rChannel_rAddr_valid,
  output [14:0]  io_mem_rChannel_rAddr_bits,
  output         io_mem_rChannel_rData_ready,
  input          io_mem_rChannel_rData_valid,
  input  [15:0]  io_mem_rChannel_rData_bits,
  input          io_mem_rChannel_rLast,
  input          io_mem_wChannel_wAddr_ready,
  output         io_mem_wChannel_wAddr_valid,
  output [14:0]  io_mem_wChannel_wAddr_bits,
  input          io_mem_wChannel_wData_ready,
  output         io_mem_wChannel_wData_valid,
  output [15:0]  io_mem_wChannel_wData_bits,
  output         io_mem_wChannel_wLast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [127:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [127:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
`endif // RANDOMIZE_REG_INIT
  wire  missQueue_clock; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_reset; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_push; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_pushEntry_rw; // @[SharedPipelinedCache.scala 49:25]
  wire [1:0] missQueue_io_pushEntry_reqId; // @[SharedPipelinedCache.scala 49:25]
  wire [1:0] missQueue_io_pushEntry_coreId; // @[SharedPipelinedCache.scala 49:25]
  wire [127:0] missQueue_io_pushEntry_wData; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_pushEntry_replaceWay; // @[SharedPipelinedCache.scala 49:25]
  wire [3:0] missQueue_io_pushEntry_tag; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_pushEntry_index; // @[SharedPipelinedCache.scala 49:25]
  wire [1:0] missQueue_io_pushEntry_blockOffset; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_pop; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_popEntry_rw; // @[SharedPipelinedCache.scala 49:25]
  wire [1:0] missQueue_io_popEntry_reqId; // @[SharedPipelinedCache.scala 49:25]
  wire [1:0] missQueue_io_popEntry_coreId; // @[SharedPipelinedCache.scala 49:25]
  wire [127:0] missQueue_io_popEntry_wData; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_popEntry_replaceWay; // @[SharedPipelinedCache.scala 49:25]
  wire [3:0] missQueue_io_popEntry_tag; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_popEntry_index; // @[SharedPipelinedCache.scala 49:25]
  wire [1:0] missQueue_io_popEntry_blockOffset; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_0; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_1; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_2; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_3; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_4; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_5; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_6; // @[SharedPipelinedCache.scala 49:25]
  wire [4:0] missQueue_io_currentIndexes_7; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_0; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_1; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_2; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_3; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_4; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_5; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_6; // @[SharedPipelinedCache.scala 49:25]
  wire [2:0] missQueue_io_currentWays_7; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_0; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_1; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_2; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_3; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_4; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_5; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_6; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_validMSHRs_7; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_full; // @[SharedPipelinedCache.scala 49:25]
  wire  missQueue_io_empty; // @[SharedPipelinedCache.scala 49:25]
  wire  updateLogic_io_readStage_valid; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_readStage_reqId; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_readStage_coreId; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_readStage_rw; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_readStage_wData; // @[SharedPipelinedCache.scala 50:27]
  wire [2:0] updateLogic_io_readStage_wWay; // @[SharedPipelinedCache.scala 50:27]
  wire [3:0] updateLogic_io_readStage_tag; // @[SharedPipelinedCache.scala 50:27]
  wire [4:0] updateLogic_io_readStage_index; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_readStage_blockOffset; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_readStage_memReadData_0; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_readStage_memReadData_1; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_readStage_memReadData_2; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_readStage_memReadData_3; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_memoryInterface_valid; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_memoryInterface_reqId; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_memoryInterface_coreId; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_memoryInterface_rw; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_memoryInterface_wData; // @[SharedPipelinedCache.scala 50:27]
  wire [2:0] updateLogic_io_memoryInterface_wWay; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_memoryInterface_responseStatus; // @[SharedPipelinedCache.scala 50:27]
  wire [3:0] updateLogic_io_memoryInterface_tag; // @[SharedPipelinedCache.scala 50:27]
  wire [4:0] updateLogic_io_memoryInterface_index; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_memoryInterface_blockOffset; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_memoryInterface_memReadData_0; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_memoryInterface_memReadData_1; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_memoryInterface_memReadData_2; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_memoryInterface_memReadData_3; // @[SharedPipelinedCache.scala 50:27]
  wire [3:0] updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 50:27]
  wire [2:0] updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_cacheUpdateControl_coreId; // @[SharedPipelinedCache.scala 50:27]
  wire [2:0] updateLogic_io_cacheUpdateControl_way; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_cacheUpdateControl_refill; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_cacheUpdateControl_update; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_cacheUpdateControl_stall; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_cacheUpdateControl_memWriteData_0; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_cacheUpdateControl_memWriteData_1; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_cacheUpdateControl_memWriteData_2; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_cacheUpdateControl_memWriteData_3; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_cacheUpdateControl_wrEn; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_coreResp_reqId_valid; // @[SharedPipelinedCache.scala 50:27]
  wire [1:0] updateLogic_io_coreResp_reqId_bits; // @[SharedPipelinedCache.scala 50:27]
  wire [127:0] updateLogic_io_coreResp_rData; // @[SharedPipelinedCache.scala 50:27]
  wire  updateLogic_io_coreResp_responseStatus; // @[SharedPipelinedCache.scala 50:27]
  wire  arbiter_clock; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_0_reqId_ready; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_0_reqId_valid; // @[SharedPipelinedCache.scala 55:23]
  wire [1:0] arbiter_io_ports_0_reqId_bits; // @[SharedPipelinedCache.scala 55:23]
  wire [14:0] arbiter_io_ports_0_addr; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_0_rw; // @[SharedPipelinedCache.scala 55:23]
  wire [127:0] arbiter_io_ports_0_wData; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_1_reqId_ready; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_1_reqId_valid; // @[SharedPipelinedCache.scala 55:23]
  wire [1:0] arbiter_io_ports_1_reqId_bits; // @[SharedPipelinedCache.scala 55:23]
  wire [14:0] arbiter_io_ports_1_addr; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_1_rw; // @[SharedPipelinedCache.scala 55:23]
  wire [127:0] arbiter_io_ports_1_wData; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_2_reqId_ready; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_2_reqId_valid; // @[SharedPipelinedCache.scala 55:23]
  wire [1:0] arbiter_io_ports_2_reqId_bits; // @[SharedPipelinedCache.scala 55:23]
  wire [14:0] arbiter_io_ports_2_addr; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_2_rw; // @[SharedPipelinedCache.scala 55:23]
  wire [127:0] arbiter_io_ports_2_wData; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_3_reqId_ready; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_3_reqId_valid; // @[SharedPipelinedCache.scala 55:23]
  wire [1:0] arbiter_io_ports_3_reqId_bits; // @[SharedPipelinedCache.scala 55:23]
  wire [14:0] arbiter_io_ports_3_addr; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_ports_3_rw; // @[SharedPipelinedCache.scala 55:23]
  wire [127:0] arbiter_io_ports_3_wData; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_out_reqId_ready; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_out_reqId_valid; // @[SharedPipelinedCache.scala 55:23]
  wire [1:0] arbiter_io_out_reqId_bits; // @[SharedPipelinedCache.scala 55:23]
  wire [14:0] arbiter_io_out_addr; // @[SharedPipelinedCache.scala 55:23]
  wire  arbiter_io_out_rw; // @[SharedPipelinedCache.scala 55:23]
  wire [127:0] arbiter_io_out_wData; // @[SharedPipelinedCache.scala 55:23]
  wire [1:0] arbiter_io_chosen; // @[SharedPipelinedCache.scala 55:23]
  wire  MemBlock_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_1_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_1_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_1_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_1_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_1_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_1_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_2_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_2_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_2_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_2_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_2_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_2_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_3_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_3_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_3_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_3_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_3_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_3_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_4_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_4_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_4_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_4_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_4_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_4_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_5_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_5_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_5_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_5_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_5_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_5_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_6_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_6_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_6_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_6_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_6_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_6_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_7_clock; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_7_io_readAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [4:0] MemBlock_7_io_writeAddr; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_7_io_writeData; // @[SharedPipelinedCache.scala 72:40]
  wire  MemBlock_7_io_wrEn; // @[SharedPipelinedCache.scala 72:40]
  wire [3:0] MemBlock_7_io_readData; // @[SharedPipelinedCache.scala 72:40]
  wire  dataMem_clock; // @[SharedPipelinedCache.scala 194:23]
  wire [4:0] dataMem_io_rIndex; // @[SharedPipelinedCache.scala 194:23]
  wire [2:0] dataMem_io_rWayIdx; // @[SharedPipelinedCache.scala 194:23]
  wire [4:0] dataMem_io_wrIndex; // @[SharedPipelinedCache.scala 194:23]
  wire [2:0] dataMem_io_wrWayIdx; // @[SharedPipelinedCache.scala 194:23]
  wire  dataMem_io_wrEn; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_wrData_0; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_wrData_1; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_wrData_2; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_wrData_3; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_rData_0; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_rData_1; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_rData_2; // @[SharedPipelinedCache.scala 194:23]
  wire [127:0] dataMem_io_rData_3; // @[SharedPipelinedCache.scala 194:23]
  wire  wbQueue_clock; // @[SharedPipelinedCache.scala 219:23]
  wire  wbQueue_reset; // @[SharedPipelinedCache.scala 219:23]
  wire  wbQueue_io_push; // @[SharedPipelinedCache.scala 219:23]
  wire  wbQueue_io_pop; // @[SharedPipelinedCache.scala 219:23]
  wire [3:0] wbQueue_io_pushEntry_tag; // @[SharedPipelinedCache.scala 219:23]
  wire [4:0] wbQueue_io_pushEntry_index; // @[SharedPipelinedCache.scala 219:23]
  wire [511:0] wbQueue_io_pushEntry_wbData; // @[SharedPipelinedCache.scala 219:23]
  wire [3:0] wbQueue_io_popEntry_tag; // @[SharedPipelinedCache.scala 219:23]
  wire [4:0] wbQueue_io_popEntry_index; // @[SharedPipelinedCache.scala 219:23]
  wire [511:0] wbQueue_io_popEntry_wbData; // @[SharedPipelinedCache.scala 219:23]
  wire  wbQueue_io_empty; // @[SharedPipelinedCache.scala 219:23]
  wire  memInterface_clock; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_reset; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_missFifo_popEntry_rw; // @[SharedPipelinedCache.scala 228:28]
  wire [1:0] memInterface_io_missFifo_popEntry_reqId; // @[SharedPipelinedCache.scala 228:28]
  wire [1:0] memInterface_io_missFifo_popEntry_coreId; // @[SharedPipelinedCache.scala 228:28]
  wire [127:0] memInterface_io_missFifo_popEntry_wData; // @[SharedPipelinedCache.scala 228:28]
  wire [2:0] memInterface_io_missFifo_popEntry_replaceWay; // @[SharedPipelinedCache.scala 228:28]
  wire [3:0] memInterface_io_missFifo_popEntry_tag; // @[SharedPipelinedCache.scala 228:28]
  wire [4:0] memInterface_io_missFifo_popEntry_index; // @[SharedPipelinedCache.scala 228:28]
  wire [1:0] memInterface_io_missFifo_popEntry_blockOffset; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_missFifo_empty; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_missFifo_pop; // @[SharedPipelinedCache.scala 228:28]
  wire [3:0] memInterface_io_wbFifo_popEntry_tag; // @[SharedPipelinedCache.scala 228:28]
  wire [4:0] memInterface_io_wbFifo_popEntry_index; // @[SharedPipelinedCache.scala 228:28]
  wire [511:0] memInterface_io_wbFifo_popEntry_wbData; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_wbFifo_empty; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_wbFifo_pop; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_updateLogic_valid; // @[SharedPipelinedCache.scala 228:28]
  wire [1:0] memInterface_io_updateLogic_reqId; // @[SharedPipelinedCache.scala 228:28]
  wire [1:0] memInterface_io_updateLogic_coreId; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_updateLogic_rw; // @[SharedPipelinedCache.scala 228:28]
  wire [127:0] memInterface_io_updateLogic_wData; // @[SharedPipelinedCache.scala 228:28]
  wire [2:0] memInterface_io_updateLogic_wWay; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_updateLogic_responseStatus; // @[SharedPipelinedCache.scala 228:28]
  wire [3:0] memInterface_io_updateLogic_tag; // @[SharedPipelinedCache.scala 228:28]
  wire [4:0] memInterface_io_updateLogic_index; // @[SharedPipelinedCache.scala 228:28]
  wire [1:0] memInterface_io_updateLogic_blockOffset; // @[SharedPipelinedCache.scala 228:28]
  wire [127:0] memInterface_io_updateLogic_memReadData_0; // @[SharedPipelinedCache.scala 228:28]
  wire [127:0] memInterface_io_updateLogic_memReadData_1; // @[SharedPipelinedCache.scala 228:28]
  wire [127:0] memInterface_io_updateLogic_memReadData_2; // @[SharedPipelinedCache.scala 228:28]
  wire [127:0] memInterface_io_updateLogic_memReadData_3; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_rChannel_rAddr_ready; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_rChannel_rAddr_valid; // @[SharedPipelinedCache.scala 228:28]
  wire [14:0] memInterface_io_memController_rChannel_rAddr_bits; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_rChannel_rData_ready; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_rChannel_rData_valid; // @[SharedPipelinedCache.scala 228:28]
  wire [15:0] memInterface_io_memController_rChannel_rData_bits; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_rChannel_rLast; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_wChannel_wAddr_ready; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_wChannel_wAddr_valid; // @[SharedPipelinedCache.scala 228:28]
  wire [14:0] memInterface_io_memController_wChannel_wAddr_bits; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_wChannel_wData_ready; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_wChannel_wData_valid; // @[SharedPipelinedCache.scala 228:28]
  wire [15:0] memInterface_io_memController_wChannel_wData_bits; // @[SharedPipelinedCache.scala 228:28]
  wire  memInterface_io_memController_wChannel_wLast; // @[SharedPipelinedCache.scala 228:28]
  wire  _reqAccept_T = ~updateLogic_io_cacheUpdateControl_stall; // @[SharedPipelinedCache.scala 56:19]
  wire  reqAccept = ~updateLogic_io_cacheUpdateControl_stall & ~missQueue_io_full; // @[SharedPipelinedCache.scala 56:30]
  wire [1:0] blockOffset = arbiter_io_out_addr[5:4]; // @[SharedPipelinedCache.scala 68:40]
  wire [4:0] index = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  wire [3:0] tag = arbiter_io_out_addr[14:11]; // @[SharedPipelinedCache.scala 70:32]
  wire  isUpdateWay = updateLogic_io_cacheUpdateControl_way == 3'h0; // @[SharedPipelinedCache.scala 76:61]
  wire  _T = updateLogic_io_cacheUpdateControl_refill & isUpdateWay; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_1 = updateLogic_io_cacheUpdateControl_way == 3'h1; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_1 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_1; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_2 = updateLogic_io_cacheUpdateControl_way == 3'h2; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_2 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_2; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_3 = updateLogic_io_cacheUpdateControl_way == 3'h3; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_3 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_3; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_4 = updateLogic_io_cacheUpdateControl_way == 3'h4; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_4 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_4; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_5 = updateLogic_io_cacheUpdateControl_way == 3'h5; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_5 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_5; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_6 = updateLogic_io_cacheUpdateControl_way == 3'h6; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_6 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_6; // @[SharedPipelinedCache.scala 82:72]
  wire  isUpdateWay_7 = updateLogic_io_cacheUpdateControl_way == 3'h7; // @[SharedPipelinedCache.scala 76:61]
  wire  _T_7 = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_7; // @[SharedPipelinedCache.scala 82:72]
  reg [1:0] coreIdTagReg; // @[SharedPipelinedCache.scala 42:30]
  wire  _reqValidTagReg_T = arbiter_io_out_reqId_valid & reqAccept; // @[SharedPipelinedCache.scala 88:63]
  reg  reqValidTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg [1:0] reqIdTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg  reqRwTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg [127:0] wDataTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg [1:0] blockTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg [4:0] indexTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] tagTagReg; // @[SharedPipelinedCache.scala 42:30]
  reg  REG__0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG__31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_1_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_2_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_3_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_4_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_5_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_6_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_0; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_1; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_2; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_3; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_4; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_5; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_6; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_7; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_8; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_9; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_10; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_11; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_12; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_13; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_14; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_15; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_16; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_17; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_18; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_19; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_20; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_21; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_22; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_23; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_24; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_25; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_26; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_27; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_28; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_29; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_30; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_7_31; // @[SharedPipelinedCache.scala 98:44]
  reg  REG_8_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_8_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_9_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_10_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_11_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_12_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_13_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_14_31; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_0; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_1; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_2; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_3; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_4; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_5; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_6; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_7; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_8; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_9; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_10; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_11; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_12; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_13; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_14; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_15; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_16; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_17; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_18; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_19; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_20; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_21; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_22; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_23; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_24; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_25; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_26; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_27; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_28; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_29; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_30; // @[SharedPipelinedCache.scala 99:44]
  reg  REG_15_31; // @[SharedPipelinedCache.scala 99:44]
  wire [3:0] readTags_0 = MemBlock_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_9 = 5'h1 == indexTagReg ? REG_8_1 : REG_8_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_10 = 5'h2 == indexTagReg ? REG_8_2 : _GEN_9; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_11 = 5'h3 == indexTagReg ? REG_8_3 : _GEN_10; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_12 = 5'h4 == indexTagReg ? REG_8_4 : _GEN_11; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_13 = 5'h5 == indexTagReg ? REG_8_5 : _GEN_12; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_14 = 5'h6 == indexTagReg ? REG_8_6 : _GEN_13; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_15 = 5'h7 == indexTagReg ? REG_8_7 : _GEN_14; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_16 = 5'h8 == indexTagReg ? REG_8_8 : _GEN_15; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_17 = 5'h9 == indexTagReg ? REG_8_9 : _GEN_16; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_18 = 5'ha == indexTagReg ? REG_8_10 : _GEN_17; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_19 = 5'hb == indexTagReg ? REG_8_11 : _GEN_18; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_20 = 5'hc == indexTagReg ? REG_8_12 : _GEN_19; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_21 = 5'hd == indexTagReg ? REG_8_13 : _GEN_20; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_22 = 5'he == indexTagReg ? REG_8_14 : _GEN_21; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_23 = 5'hf == indexTagReg ? REG_8_15 : _GEN_22; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_24 = 5'h10 == indexTagReg ? REG_8_16 : _GEN_23; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_25 = 5'h11 == indexTagReg ? REG_8_17 : _GEN_24; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_26 = 5'h12 == indexTagReg ? REG_8_18 : _GEN_25; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_27 = 5'h13 == indexTagReg ? REG_8_19 : _GEN_26; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_28 = 5'h14 == indexTagReg ? REG_8_20 : _GEN_27; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_29 = 5'h15 == indexTagReg ? REG_8_21 : _GEN_28; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_30 = 5'h16 == indexTagReg ? REG_8_22 : _GEN_29; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_31 = 5'h17 == indexTagReg ? REG_8_23 : _GEN_30; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_32 = 5'h18 == indexTagReg ? REG_8_24 : _GEN_31; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_33 = 5'h19 == indexTagReg ? REG_8_25 : _GEN_32; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_34 = 5'h1a == indexTagReg ? REG_8_26 : _GEN_33; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_35 = 5'h1b == indexTagReg ? REG_8_27 : _GEN_34; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_36 = 5'h1c == indexTagReg ? REG_8_28 : _GEN_35; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_37 = 5'h1d == indexTagReg ? REG_8_29 : _GEN_36; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_38 = 5'h1e == indexTagReg ? REG_8_30 : _GEN_37; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_39 = 5'h1f == indexTagReg ? REG_8_31 : _GEN_38; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_0 = _GEN_39 & tagTagReg == readTags_0; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_41 = 5'h1 == indexTagReg ? REG__1 : REG__0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_42 = 5'h2 == indexTagReg ? REG__2 : _GEN_41; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_43 = 5'h3 == indexTagReg ? REG__3 : _GEN_42; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_44 = 5'h4 == indexTagReg ? REG__4 : _GEN_43; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_45 = 5'h5 == indexTagReg ? REG__5 : _GEN_44; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_46 = 5'h6 == indexTagReg ? REG__6 : _GEN_45; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_47 = 5'h7 == indexTagReg ? REG__7 : _GEN_46; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_48 = 5'h8 == indexTagReg ? REG__8 : _GEN_47; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_49 = 5'h9 == indexTagReg ? REG__9 : _GEN_48; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_50 = 5'ha == indexTagReg ? REG__10 : _GEN_49; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_51 = 5'hb == indexTagReg ? REG__11 : _GEN_50; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_52 = 5'hc == indexTagReg ? REG__12 : _GEN_51; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_53 = 5'hd == indexTagReg ? REG__13 : _GEN_52; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_54 = 5'he == indexTagReg ? REG__14 : _GEN_53; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_55 = 5'hf == indexTagReg ? REG__15 : _GEN_54; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_56 = 5'h10 == indexTagReg ? REG__16 : _GEN_55; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_57 = 5'h11 == indexTagReg ? REG__17 : _GEN_56; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_58 = 5'h12 == indexTagReg ? REG__18 : _GEN_57; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_59 = 5'h13 == indexTagReg ? REG__19 : _GEN_58; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_60 = 5'h14 == indexTagReg ? REG__20 : _GEN_59; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_61 = 5'h15 == indexTagReg ? REG__21 : _GEN_60; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_62 = 5'h16 == indexTagReg ? REG__22 : _GEN_61; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_63 = 5'h17 == indexTagReg ? REG__23 : _GEN_62; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_64 = 5'h18 == indexTagReg ? REG__24 : _GEN_63; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_65 = 5'h19 == indexTagReg ? REG__25 : _GEN_64; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_66 = 5'h1a == indexTagReg ? REG__26 : _GEN_65; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_67 = 5'h1b == indexTagReg ? REG__27 : _GEN_66; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_68 = 5'h1c == indexTagReg ? REG__28 : _GEN_67; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_69 = 5'h1d == indexTagReg ? REG__29 : _GEN_68; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2624 = 3'h0 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_72 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_8_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2625 = 3'h1 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_73 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_8_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2626 = 3'h2 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_74 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_8_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2627 = 3'h3 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_75 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_8_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2628 = 3'h4 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_76 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_8_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2629 = 3'h5 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_77 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_8_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2630 = 3'h6 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_78 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_8_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2631 = 3'h7 == updateLogic_io_cacheUpdateControl_index; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_79 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_8_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire [3:0] _GEN_2632 = {{1'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2633 = 4'h8 == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_80 = 4'h8 == _GEN_2632 | REG_8_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2635 = 4'h9 == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_81 = 4'h9 == _GEN_2632 | REG_8_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2637 = 4'ha == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_82 = 4'ha == _GEN_2632 | REG_8_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2639 = 4'hb == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_83 = 4'hb == _GEN_2632 | REG_8_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2641 = 4'hc == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_84 = 4'hc == _GEN_2632 | REG_8_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2643 = 4'hd == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_85 = 4'hd == _GEN_2632 | REG_8_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2645 = 4'he == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_86 = 4'he == _GEN_2632 | REG_8_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2647 = 4'hf == _GEN_2632; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_87 = 4'hf == _GEN_2632 | REG_8_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire [4:0] _GEN_2648 = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2649 = 5'h10 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_88 = 5'h10 == _GEN_2648 | REG_8_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2651 = 5'h11 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_89 = 5'h11 == _GEN_2648 | REG_8_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2653 = 5'h12 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_90 = 5'h12 == _GEN_2648 | REG_8_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2655 = 5'h13 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_91 = 5'h13 == _GEN_2648 | REG_8_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2657 = 5'h14 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_92 = 5'h14 == _GEN_2648 | REG_8_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2659 = 5'h15 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_93 = 5'h15 == _GEN_2648 | REG_8_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2661 = 5'h16 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_94 = 5'h16 == _GEN_2648 | REG_8_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2663 = 5'h17 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_95 = 5'h17 == _GEN_2648 | REG_8_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2665 = 5'h18 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_96 = 5'h18 == _GEN_2648 | REG_8_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2667 = 5'h19 == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_97 = 5'h19 == _GEN_2648 | REG_8_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2669 = 5'h1a == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_98 = 5'h1a == _GEN_2648 | REG_8_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2671 = 5'h1b == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_99 = 5'h1b == _GEN_2648 | REG_8_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2673 = 5'h1c == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_100 = 5'h1c == _GEN_2648 | REG_8_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2675 = 5'h1d == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_101 = 5'h1d == _GEN_2648 | REG_8_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2677 = 5'h1e == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_102 = 5'h1e == _GEN_2648 | REG_8_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2679 = 5'h1f == _GEN_2648; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_103 = 5'h1f == _GEN_2648 | REG_8_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_104 = _GEN_2624 | REG__0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_105 = _GEN_2625 | REG__1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_106 = _GEN_2626 | REG__2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_107 = _GEN_2627 | REG__3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_108 = _GEN_2628 | REG__4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_109 = _GEN_2629 | REG__5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_110 = _GEN_2630 | REG__6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_111 = _GEN_2631 | REG__7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_112 = _GEN_2633 | REG__8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_113 = _GEN_2635 | REG__9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_114 = _GEN_2637 | REG__10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_115 = _GEN_2639 | REG__11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_116 = _GEN_2641 | REG__12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_117 = _GEN_2643 | REG__13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_118 = _GEN_2645 | REG__14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_119 = _GEN_2647 | REG__15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_120 = _GEN_2649 | REG__16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_121 = _GEN_2651 | REG__17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_122 = _GEN_2653 | REG__18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_123 = _GEN_2655 | REG__19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_124 = _GEN_2657 | REG__20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_125 = _GEN_2659 | REG__21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_126 = _GEN_2661 | REG__22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_127 = _GEN_2663 | REG__23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_128 = _GEN_2665 | REG__24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_129 = _GEN_2667 | REG__25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_130 = _GEN_2669 | REG__26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_131 = _GEN_2671 | REG__27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_132 = _GEN_2673 | REG__28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_133 = _GEN_2675 | REG__29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_134 = _GEN_2677 | REG__30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_135 = _GEN_2679 | REG__31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_136 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_137 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_138 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_139 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_140 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_141 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_142 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_143 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG__7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_144 = 4'h8 == _GEN_2632 ? 1'h0 : REG__8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_145 = 4'h9 == _GEN_2632 ? 1'h0 : REG__9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_146 = 4'ha == _GEN_2632 ? 1'h0 : REG__10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_147 = 4'hb == _GEN_2632 ? 1'h0 : REG__11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_148 = 4'hc == _GEN_2632 ? 1'h0 : REG__12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_149 = 4'hd == _GEN_2632 ? 1'h0 : REG__13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_150 = 4'he == _GEN_2632 ? 1'h0 : REG__14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_151 = 4'hf == _GEN_2632 ? 1'h0 : REG__15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_152 = 5'h10 == _GEN_2648 ? 1'h0 : REG__16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_153 = 5'h11 == _GEN_2648 ? 1'h0 : REG__17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_154 = 5'h12 == _GEN_2648 ? 1'h0 : REG__18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_155 = 5'h13 == _GEN_2648 ? 1'h0 : REG__19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_156 = 5'h14 == _GEN_2648 ? 1'h0 : REG__20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_157 = 5'h15 == _GEN_2648 ? 1'h0 : REG__21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_158 = 5'h16 == _GEN_2648 ? 1'h0 : REG__22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_159 = 5'h17 == _GEN_2648 ? 1'h0 : REG__23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_160 = 5'h18 == _GEN_2648 ? 1'h0 : REG__24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_161 = 5'h19 == _GEN_2648 ? 1'h0 : REG__25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_162 = 5'h1a == _GEN_2648 ? 1'h0 : REG__26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_163 = 5'h1b == _GEN_2648 ? 1'h0 : REG__27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_164 = 5'h1c == _GEN_2648 ? 1'h0 : REG__28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_165 = 5'h1d == _GEN_2648 ? 1'h0 : REG__29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_166 = 5'h1e == _GEN_2648 ? 1'h0 : REG__30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_167 = 5'h1f == _GEN_2648 ? 1'h0 : REG__31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_168 = updateLogic_io_cacheUpdateControl_update ? _GEN_104 : _GEN_136; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_169 = updateLogic_io_cacheUpdateControl_update ? _GEN_105 : _GEN_137; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_170 = updateLogic_io_cacheUpdateControl_update ? _GEN_106 : _GEN_138; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_171 = updateLogic_io_cacheUpdateControl_update ? _GEN_107 : _GEN_139; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_172 = updateLogic_io_cacheUpdateControl_update ? _GEN_108 : _GEN_140; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_173 = updateLogic_io_cacheUpdateControl_update ? _GEN_109 : _GEN_141; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_174 = updateLogic_io_cacheUpdateControl_update ? _GEN_110 : _GEN_142; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_175 = updateLogic_io_cacheUpdateControl_update ? _GEN_111 : _GEN_143; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_176 = updateLogic_io_cacheUpdateControl_update ? _GEN_112 : _GEN_144; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_177 = updateLogic_io_cacheUpdateControl_update ? _GEN_113 : _GEN_145; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_178 = updateLogic_io_cacheUpdateControl_update ? _GEN_114 : _GEN_146; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_179 = updateLogic_io_cacheUpdateControl_update ? _GEN_115 : _GEN_147; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_180 = updateLogic_io_cacheUpdateControl_update ? _GEN_116 : _GEN_148; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_181 = updateLogic_io_cacheUpdateControl_update ? _GEN_117 : _GEN_149; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_182 = updateLogic_io_cacheUpdateControl_update ? _GEN_118 : _GEN_150; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_183 = updateLogic_io_cacheUpdateControl_update ? _GEN_119 : _GEN_151; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_184 = updateLogic_io_cacheUpdateControl_update ? _GEN_120 : _GEN_152; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_185 = updateLogic_io_cacheUpdateControl_update ? _GEN_121 : _GEN_153; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_186 = updateLogic_io_cacheUpdateControl_update ? _GEN_122 : _GEN_154; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_187 = updateLogic_io_cacheUpdateControl_update ? _GEN_123 : _GEN_155; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_188 = updateLogic_io_cacheUpdateControl_update ? _GEN_124 : _GEN_156; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_189 = updateLogic_io_cacheUpdateControl_update ? _GEN_125 : _GEN_157; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_190 = updateLogic_io_cacheUpdateControl_update ? _GEN_126 : _GEN_158; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_191 = updateLogic_io_cacheUpdateControl_update ? _GEN_127 : _GEN_159; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_192 = updateLogic_io_cacheUpdateControl_update ? _GEN_128 : _GEN_160; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_193 = updateLogic_io_cacheUpdateControl_update ? _GEN_129 : _GEN_161; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_194 = updateLogic_io_cacheUpdateControl_update ? _GEN_130 : _GEN_162; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_195 = updateLogic_io_cacheUpdateControl_update ? _GEN_131 : _GEN_163; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_196 = updateLogic_io_cacheUpdateControl_update ? _GEN_132 : _GEN_164; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_197 = updateLogic_io_cacheUpdateControl_update ? _GEN_133 : _GEN_165; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_198 = updateLogic_io_cacheUpdateControl_update ? _GEN_134 : _GEN_166; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_199 = updateLogic_io_cacheUpdateControl_update ? _GEN_135 : _GEN_167; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_232 = _T ? _GEN_168 : REG__0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_233 = _T ? _GEN_169 : REG__1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_234 = _T ? _GEN_170 : REG__2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_235 = _T ? _GEN_171 : REG__3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_236 = _T ? _GEN_172 : REG__4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_237 = _T ? _GEN_173 : REG__5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_238 = _T ? _GEN_174 : REG__6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_239 = _T ? _GEN_175 : REG__7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_240 = _T ? _GEN_176 : REG__8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_241 = _T ? _GEN_177 : REG__9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_242 = _T ? _GEN_178 : REG__10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_243 = _T ? _GEN_179 : REG__11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_244 = _T ? _GEN_180 : REG__12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_245 = _T ? _GEN_181 : REG__13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_246 = _T ? _GEN_182 : REG__14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_247 = _T ? _GEN_183 : REG__15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_248 = _T ? _GEN_184 : REG__16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_249 = _T ? _GEN_185 : REG__17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_250 = _T ? _GEN_186 : REG__18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_251 = _T ? _GEN_187 : REG__19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_252 = _T ? _GEN_188 : REG__20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_253 = _T ? _GEN_189 : REG__21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_254 = _T ? _GEN_190 : REG__22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_255 = _T ? _GEN_191 : REG__23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_256 = _T ? _GEN_192 : REG__24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_257 = _T ? _GEN_193 : REG__25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_258 = _T ? _GEN_194 : REG__26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_259 = _T ? _GEN_195 : REG__27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_260 = _T ? _GEN_196 : REG__28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_261 = _T ? _GEN_197 : REG__29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_262 = _T ? _GEN_198 : REG__30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_263 = _T ? _GEN_199 : REG__31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_264 = _GEN_2624 | _GEN_232; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_265 = _GEN_2625 | _GEN_233; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_266 = _GEN_2626 | _GEN_234; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_267 = _GEN_2627 | _GEN_235; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_268 = _GEN_2628 | _GEN_236; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_269 = _GEN_2629 | _GEN_237; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_270 = _GEN_2630 | _GEN_238; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_271 = _GEN_2631 | _GEN_239; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_272 = _GEN_2633 | _GEN_240; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_273 = _GEN_2635 | _GEN_241; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_274 = _GEN_2637 | _GEN_242; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_275 = _GEN_2639 | _GEN_243; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_276 = _GEN_2641 | _GEN_244; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_277 = _GEN_2643 | _GEN_245; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_278 = _GEN_2645 | _GEN_246; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_279 = _GEN_2647 | _GEN_247; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_280 = _GEN_2649 | _GEN_248; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_281 = _GEN_2651 | _GEN_249; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_282 = _GEN_2653 | _GEN_250; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_283 = _GEN_2655 | _GEN_251; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_284 = _GEN_2657 | _GEN_252; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_285 = _GEN_2659 | _GEN_253; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_286 = _GEN_2661 | _GEN_254; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_287 = _GEN_2663 | _GEN_255; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_288 = _GEN_2665 | _GEN_256; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_289 = _GEN_2667 | _GEN_257; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_290 = _GEN_2669 | _GEN_258; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_291 = _GEN_2671 | _GEN_259; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_292 = _GEN_2673 | _GEN_260; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_293 = _GEN_2675 | _GEN_261; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_294 = _GEN_2677 | _GEN_262; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_295 = _GEN_2679 | _GEN_263; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_1 = MemBlock_1_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_329 = 5'h1 == indexTagReg ? REG_9_1 : REG_9_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_330 = 5'h2 == indexTagReg ? REG_9_2 : _GEN_329; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_331 = 5'h3 == indexTagReg ? REG_9_3 : _GEN_330; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_332 = 5'h4 == indexTagReg ? REG_9_4 : _GEN_331; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_333 = 5'h5 == indexTagReg ? REG_9_5 : _GEN_332; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_334 = 5'h6 == indexTagReg ? REG_9_6 : _GEN_333; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_335 = 5'h7 == indexTagReg ? REG_9_7 : _GEN_334; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_336 = 5'h8 == indexTagReg ? REG_9_8 : _GEN_335; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_337 = 5'h9 == indexTagReg ? REG_9_9 : _GEN_336; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_338 = 5'ha == indexTagReg ? REG_9_10 : _GEN_337; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_339 = 5'hb == indexTagReg ? REG_9_11 : _GEN_338; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_340 = 5'hc == indexTagReg ? REG_9_12 : _GEN_339; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_341 = 5'hd == indexTagReg ? REG_9_13 : _GEN_340; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_342 = 5'he == indexTagReg ? REG_9_14 : _GEN_341; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_343 = 5'hf == indexTagReg ? REG_9_15 : _GEN_342; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_344 = 5'h10 == indexTagReg ? REG_9_16 : _GEN_343; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_345 = 5'h11 == indexTagReg ? REG_9_17 : _GEN_344; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_346 = 5'h12 == indexTagReg ? REG_9_18 : _GEN_345; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_347 = 5'h13 == indexTagReg ? REG_9_19 : _GEN_346; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_348 = 5'h14 == indexTagReg ? REG_9_20 : _GEN_347; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_349 = 5'h15 == indexTagReg ? REG_9_21 : _GEN_348; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_350 = 5'h16 == indexTagReg ? REG_9_22 : _GEN_349; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_351 = 5'h17 == indexTagReg ? REG_9_23 : _GEN_350; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_352 = 5'h18 == indexTagReg ? REG_9_24 : _GEN_351; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_353 = 5'h19 == indexTagReg ? REG_9_25 : _GEN_352; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_354 = 5'h1a == indexTagReg ? REG_9_26 : _GEN_353; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_355 = 5'h1b == indexTagReg ? REG_9_27 : _GEN_354; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_356 = 5'h1c == indexTagReg ? REG_9_28 : _GEN_355; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_357 = 5'h1d == indexTagReg ? REG_9_29 : _GEN_356; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_358 = 5'h1e == indexTagReg ? REG_9_30 : _GEN_357; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_359 = 5'h1f == indexTagReg ? REG_9_31 : _GEN_358; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_1 = _GEN_359 & tagTagReg == readTags_1; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_361 = 5'h1 == indexTagReg ? REG_1_1 : REG_1_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_362 = 5'h2 == indexTagReg ? REG_1_2 : _GEN_361; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_363 = 5'h3 == indexTagReg ? REG_1_3 : _GEN_362; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_364 = 5'h4 == indexTagReg ? REG_1_4 : _GEN_363; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_365 = 5'h5 == indexTagReg ? REG_1_5 : _GEN_364; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_366 = 5'h6 == indexTagReg ? REG_1_6 : _GEN_365; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_367 = 5'h7 == indexTagReg ? REG_1_7 : _GEN_366; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_368 = 5'h8 == indexTagReg ? REG_1_8 : _GEN_367; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_369 = 5'h9 == indexTagReg ? REG_1_9 : _GEN_368; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_370 = 5'ha == indexTagReg ? REG_1_10 : _GEN_369; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_371 = 5'hb == indexTagReg ? REG_1_11 : _GEN_370; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_372 = 5'hc == indexTagReg ? REG_1_12 : _GEN_371; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_373 = 5'hd == indexTagReg ? REG_1_13 : _GEN_372; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_374 = 5'he == indexTagReg ? REG_1_14 : _GEN_373; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_375 = 5'hf == indexTagReg ? REG_1_15 : _GEN_374; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_376 = 5'h10 == indexTagReg ? REG_1_16 : _GEN_375; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_377 = 5'h11 == indexTagReg ? REG_1_17 : _GEN_376; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_378 = 5'h12 == indexTagReg ? REG_1_18 : _GEN_377; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_379 = 5'h13 == indexTagReg ? REG_1_19 : _GEN_378; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_380 = 5'h14 == indexTagReg ? REG_1_20 : _GEN_379; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_381 = 5'h15 == indexTagReg ? REG_1_21 : _GEN_380; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_382 = 5'h16 == indexTagReg ? REG_1_22 : _GEN_381; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_383 = 5'h17 == indexTagReg ? REG_1_23 : _GEN_382; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_384 = 5'h18 == indexTagReg ? REG_1_24 : _GEN_383; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_385 = 5'h19 == indexTagReg ? REG_1_25 : _GEN_384; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_386 = 5'h1a == indexTagReg ? REG_1_26 : _GEN_385; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_387 = 5'h1b == indexTagReg ? REG_1_27 : _GEN_386; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_388 = 5'h1c == indexTagReg ? REG_1_28 : _GEN_387; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_389 = 5'h1d == indexTagReg ? REG_1_29 : _GEN_388; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_392 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_9_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_393 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_9_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_394 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_9_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_395 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_9_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_396 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_9_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_397 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_9_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_398 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_9_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_399 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_9_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_400 = 4'h8 == _GEN_2632 | REG_9_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_401 = 4'h9 == _GEN_2632 | REG_9_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_402 = 4'ha == _GEN_2632 | REG_9_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_403 = 4'hb == _GEN_2632 | REG_9_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_404 = 4'hc == _GEN_2632 | REG_9_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_405 = 4'hd == _GEN_2632 | REG_9_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_406 = 4'he == _GEN_2632 | REG_9_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_407 = 4'hf == _GEN_2632 | REG_9_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_408 = 5'h10 == _GEN_2648 | REG_9_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_409 = 5'h11 == _GEN_2648 | REG_9_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_410 = 5'h12 == _GEN_2648 | REG_9_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_411 = 5'h13 == _GEN_2648 | REG_9_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_412 = 5'h14 == _GEN_2648 | REG_9_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_413 = 5'h15 == _GEN_2648 | REG_9_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_414 = 5'h16 == _GEN_2648 | REG_9_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_415 = 5'h17 == _GEN_2648 | REG_9_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_416 = 5'h18 == _GEN_2648 | REG_9_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_417 = 5'h19 == _GEN_2648 | REG_9_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_418 = 5'h1a == _GEN_2648 | REG_9_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_419 = 5'h1b == _GEN_2648 | REG_9_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_420 = 5'h1c == _GEN_2648 | REG_9_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_421 = 5'h1d == _GEN_2648 | REG_9_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_422 = 5'h1e == _GEN_2648 | REG_9_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_423 = 5'h1f == _GEN_2648 | REG_9_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_424 = _GEN_2624 | REG_1_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_425 = _GEN_2625 | REG_1_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_426 = _GEN_2626 | REG_1_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_427 = _GEN_2627 | REG_1_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_428 = _GEN_2628 | REG_1_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_429 = _GEN_2629 | REG_1_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_430 = _GEN_2630 | REG_1_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_431 = _GEN_2631 | REG_1_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_432 = _GEN_2633 | REG_1_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_433 = _GEN_2635 | REG_1_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_434 = _GEN_2637 | REG_1_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_435 = _GEN_2639 | REG_1_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_436 = _GEN_2641 | REG_1_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_437 = _GEN_2643 | REG_1_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_438 = _GEN_2645 | REG_1_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_439 = _GEN_2647 | REG_1_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_440 = _GEN_2649 | REG_1_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_441 = _GEN_2651 | REG_1_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_442 = _GEN_2653 | REG_1_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_443 = _GEN_2655 | REG_1_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_444 = _GEN_2657 | REG_1_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_445 = _GEN_2659 | REG_1_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_446 = _GEN_2661 | REG_1_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_447 = _GEN_2663 | REG_1_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_448 = _GEN_2665 | REG_1_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_449 = _GEN_2667 | REG_1_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_450 = _GEN_2669 | REG_1_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_451 = _GEN_2671 | REG_1_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_452 = _GEN_2673 | REG_1_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_453 = _GEN_2675 | REG_1_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_454 = _GEN_2677 | REG_1_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_455 = _GEN_2679 | REG_1_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_456 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_457 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_458 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_459 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_460 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_461 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_462 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_463 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_1_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_464 = 4'h8 == _GEN_2632 ? 1'h0 : REG_1_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_465 = 4'h9 == _GEN_2632 ? 1'h0 : REG_1_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_466 = 4'ha == _GEN_2632 ? 1'h0 : REG_1_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_467 = 4'hb == _GEN_2632 ? 1'h0 : REG_1_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_468 = 4'hc == _GEN_2632 ? 1'h0 : REG_1_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_469 = 4'hd == _GEN_2632 ? 1'h0 : REG_1_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_470 = 4'he == _GEN_2632 ? 1'h0 : REG_1_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_471 = 4'hf == _GEN_2632 ? 1'h0 : REG_1_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_472 = 5'h10 == _GEN_2648 ? 1'h0 : REG_1_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_473 = 5'h11 == _GEN_2648 ? 1'h0 : REG_1_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_474 = 5'h12 == _GEN_2648 ? 1'h0 : REG_1_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_475 = 5'h13 == _GEN_2648 ? 1'h0 : REG_1_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_476 = 5'h14 == _GEN_2648 ? 1'h0 : REG_1_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_477 = 5'h15 == _GEN_2648 ? 1'h0 : REG_1_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_478 = 5'h16 == _GEN_2648 ? 1'h0 : REG_1_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_479 = 5'h17 == _GEN_2648 ? 1'h0 : REG_1_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_480 = 5'h18 == _GEN_2648 ? 1'h0 : REG_1_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_481 = 5'h19 == _GEN_2648 ? 1'h0 : REG_1_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_482 = 5'h1a == _GEN_2648 ? 1'h0 : REG_1_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_483 = 5'h1b == _GEN_2648 ? 1'h0 : REG_1_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_484 = 5'h1c == _GEN_2648 ? 1'h0 : REG_1_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_485 = 5'h1d == _GEN_2648 ? 1'h0 : REG_1_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_486 = 5'h1e == _GEN_2648 ? 1'h0 : REG_1_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_487 = 5'h1f == _GEN_2648 ? 1'h0 : REG_1_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_488 = updateLogic_io_cacheUpdateControl_update ? _GEN_424 : _GEN_456; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_489 = updateLogic_io_cacheUpdateControl_update ? _GEN_425 : _GEN_457; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_490 = updateLogic_io_cacheUpdateControl_update ? _GEN_426 : _GEN_458; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_491 = updateLogic_io_cacheUpdateControl_update ? _GEN_427 : _GEN_459; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_492 = updateLogic_io_cacheUpdateControl_update ? _GEN_428 : _GEN_460; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_493 = updateLogic_io_cacheUpdateControl_update ? _GEN_429 : _GEN_461; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_494 = updateLogic_io_cacheUpdateControl_update ? _GEN_430 : _GEN_462; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_495 = updateLogic_io_cacheUpdateControl_update ? _GEN_431 : _GEN_463; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_496 = updateLogic_io_cacheUpdateControl_update ? _GEN_432 : _GEN_464; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_497 = updateLogic_io_cacheUpdateControl_update ? _GEN_433 : _GEN_465; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_498 = updateLogic_io_cacheUpdateControl_update ? _GEN_434 : _GEN_466; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_499 = updateLogic_io_cacheUpdateControl_update ? _GEN_435 : _GEN_467; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_500 = updateLogic_io_cacheUpdateControl_update ? _GEN_436 : _GEN_468; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_501 = updateLogic_io_cacheUpdateControl_update ? _GEN_437 : _GEN_469; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_502 = updateLogic_io_cacheUpdateControl_update ? _GEN_438 : _GEN_470; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_503 = updateLogic_io_cacheUpdateControl_update ? _GEN_439 : _GEN_471; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_504 = updateLogic_io_cacheUpdateControl_update ? _GEN_440 : _GEN_472; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_505 = updateLogic_io_cacheUpdateControl_update ? _GEN_441 : _GEN_473; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_506 = updateLogic_io_cacheUpdateControl_update ? _GEN_442 : _GEN_474; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_507 = updateLogic_io_cacheUpdateControl_update ? _GEN_443 : _GEN_475; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_508 = updateLogic_io_cacheUpdateControl_update ? _GEN_444 : _GEN_476; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_509 = updateLogic_io_cacheUpdateControl_update ? _GEN_445 : _GEN_477; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_510 = updateLogic_io_cacheUpdateControl_update ? _GEN_446 : _GEN_478; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_511 = updateLogic_io_cacheUpdateControl_update ? _GEN_447 : _GEN_479; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_512 = updateLogic_io_cacheUpdateControl_update ? _GEN_448 : _GEN_480; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_513 = updateLogic_io_cacheUpdateControl_update ? _GEN_449 : _GEN_481; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_514 = updateLogic_io_cacheUpdateControl_update ? _GEN_450 : _GEN_482; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_515 = updateLogic_io_cacheUpdateControl_update ? _GEN_451 : _GEN_483; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_516 = updateLogic_io_cacheUpdateControl_update ? _GEN_452 : _GEN_484; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_517 = updateLogic_io_cacheUpdateControl_update ? _GEN_453 : _GEN_485; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_518 = updateLogic_io_cacheUpdateControl_update ? _GEN_454 : _GEN_486; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_519 = updateLogic_io_cacheUpdateControl_update ? _GEN_455 : _GEN_487; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_552 = _T_1 ? _GEN_488 : REG_1_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_553 = _T_1 ? _GEN_489 : REG_1_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_554 = _T_1 ? _GEN_490 : REG_1_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_555 = _T_1 ? _GEN_491 : REG_1_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_556 = _T_1 ? _GEN_492 : REG_1_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_557 = _T_1 ? _GEN_493 : REG_1_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_558 = _T_1 ? _GEN_494 : REG_1_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_559 = _T_1 ? _GEN_495 : REG_1_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_560 = _T_1 ? _GEN_496 : REG_1_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_561 = _T_1 ? _GEN_497 : REG_1_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_562 = _T_1 ? _GEN_498 : REG_1_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_563 = _T_1 ? _GEN_499 : REG_1_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_564 = _T_1 ? _GEN_500 : REG_1_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_565 = _T_1 ? _GEN_501 : REG_1_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_566 = _T_1 ? _GEN_502 : REG_1_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_567 = _T_1 ? _GEN_503 : REG_1_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_568 = _T_1 ? _GEN_504 : REG_1_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_569 = _T_1 ? _GEN_505 : REG_1_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_570 = _T_1 ? _GEN_506 : REG_1_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_571 = _T_1 ? _GEN_507 : REG_1_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_572 = _T_1 ? _GEN_508 : REG_1_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_573 = _T_1 ? _GEN_509 : REG_1_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_574 = _T_1 ? _GEN_510 : REG_1_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_575 = _T_1 ? _GEN_511 : REG_1_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_576 = _T_1 ? _GEN_512 : REG_1_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_577 = _T_1 ? _GEN_513 : REG_1_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_578 = _T_1 ? _GEN_514 : REG_1_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_579 = _T_1 ? _GEN_515 : REG_1_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_580 = _T_1 ? _GEN_516 : REG_1_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_581 = _T_1 ? _GEN_517 : REG_1_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_582 = _T_1 ? _GEN_518 : REG_1_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_583 = _T_1 ? _GEN_519 : REG_1_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_584 = _GEN_2624 | _GEN_552; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_585 = _GEN_2625 | _GEN_553; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_586 = _GEN_2626 | _GEN_554; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_587 = _GEN_2627 | _GEN_555; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_588 = _GEN_2628 | _GEN_556; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_589 = _GEN_2629 | _GEN_557; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_590 = _GEN_2630 | _GEN_558; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_591 = _GEN_2631 | _GEN_559; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_592 = _GEN_2633 | _GEN_560; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_593 = _GEN_2635 | _GEN_561; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_594 = _GEN_2637 | _GEN_562; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_595 = _GEN_2639 | _GEN_563; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_596 = _GEN_2641 | _GEN_564; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_597 = _GEN_2643 | _GEN_565; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_598 = _GEN_2645 | _GEN_566; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_599 = _GEN_2647 | _GEN_567; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_600 = _GEN_2649 | _GEN_568; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_601 = _GEN_2651 | _GEN_569; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_602 = _GEN_2653 | _GEN_570; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_603 = _GEN_2655 | _GEN_571; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_604 = _GEN_2657 | _GEN_572; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_605 = _GEN_2659 | _GEN_573; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_606 = _GEN_2661 | _GEN_574; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_607 = _GEN_2663 | _GEN_575; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_608 = _GEN_2665 | _GEN_576; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_609 = _GEN_2667 | _GEN_577; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_610 = _GEN_2669 | _GEN_578; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_611 = _GEN_2671 | _GEN_579; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_612 = _GEN_2673 | _GEN_580; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_613 = _GEN_2675 | _GEN_581; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_614 = _GEN_2677 | _GEN_582; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_615 = _GEN_2679 | _GEN_583; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_2 = MemBlock_2_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_649 = 5'h1 == indexTagReg ? REG_10_1 : REG_10_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_650 = 5'h2 == indexTagReg ? REG_10_2 : _GEN_649; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_651 = 5'h3 == indexTagReg ? REG_10_3 : _GEN_650; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_652 = 5'h4 == indexTagReg ? REG_10_4 : _GEN_651; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_653 = 5'h5 == indexTagReg ? REG_10_5 : _GEN_652; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_654 = 5'h6 == indexTagReg ? REG_10_6 : _GEN_653; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_655 = 5'h7 == indexTagReg ? REG_10_7 : _GEN_654; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_656 = 5'h8 == indexTagReg ? REG_10_8 : _GEN_655; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_657 = 5'h9 == indexTagReg ? REG_10_9 : _GEN_656; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_658 = 5'ha == indexTagReg ? REG_10_10 : _GEN_657; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_659 = 5'hb == indexTagReg ? REG_10_11 : _GEN_658; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_660 = 5'hc == indexTagReg ? REG_10_12 : _GEN_659; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_661 = 5'hd == indexTagReg ? REG_10_13 : _GEN_660; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_662 = 5'he == indexTagReg ? REG_10_14 : _GEN_661; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_663 = 5'hf == indexTagReg ? REG_10_15 : _GEN_662; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_664 = 5'h10 == indexTagReg ? REG_10_16 : _GEN_663; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_665 = 5'h11 == indexTagReg ? REG_10_17 : _GEN_664; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_666 = 5'h12 == indexTagReg ? REG_10_18 : _GEN_665; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_667 = 5'h13 == indexTagReg ? REG_10_19 : _GEN_666; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_668 = 5'h14 == indexTagReg ? REG_10_20 : _GEN_667; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_669 = 5'h15 == indexTagReg ? REG_10_21 : _GEN_668; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_670 = 5'h16 == indexTagReg ? REG_10_22 : _GEN_669; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_671 = 5'h17 == indexTagReg ? REG_10_23 : _GEN_670; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_672 = 5'h18 == indexTagReg ? REG_10_24 : _GEN_671; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_673 = 5'h19 == indexTagReg ? REG_10_25 : _GEN_672; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_674 = 5'h1a == indexTagReg ? REG_10_26 : _GEN_673; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_675 = 5'h1b == indexTagReg ? REG_10_27 : _GEN_674; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_676 = 5'h1c == indexTagReg ? REG_10_28 : _GEN_675; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_677 = 5'h1d == indexTagReg ? REG_10_29 : _GEN_676; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_678 = 5'h1e == indexTagReg ? REG_10_30 : _GEN_677; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_679 = 5'h1f == indexTagReg ? REG_10_31 : _GEN_678; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_2 = _GEN_679 & tagTagReg == readTags_2; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_681 = 5'h1 == indexTagReg ? REG_2_1 : REG_2_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_682 = 5'h2 == indexTagReg ? REG_2_2 : _GEN_681; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_683 = 5'h3 == indexTagReg ? REG_2_3 : _GEN_682; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_684 = 5'h4 == indexTagReg ? REG_2_4 : _GEN_683; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_685 = 5'h5 == indexTagReg ? REG_2_5 : _GEN_684; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_686 = 5'h6 == indexTagReg ? REG_2_6 : _GEN_685; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_687 = 5'h7 == indexTagReg ? REG_2_7 : _GEN_686; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_688 = 5'h8 == indexTagReg ? REG_2_8 : _GEN_687; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_689 = 5'h9 == indexTagReg ? REG_2_9 : _GEN_688; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_690 = 5'ha == indexTagReg ? REG_2_10 : _GEN_689; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_691 = 5'hb == indexTagReg ? REG_2_11 : _GEN_690; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_692 = 5'hc == indexTagReg ? REG_2_12 : _GEN_691; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_693 = 5'hd == indexTagReg ? REG_2_13 : _GEN_692; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_694 = 5'he == indexTagReg ? REG_2_14 : _GEN_693; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_695 = 5'hf == indexTagReg ? REG_2_15 : _GEN_694; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_696 = 5'h10 == indexTagReg ? REG_2_16 : _GEN_695; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_697 = 5'h11 == indexTagReg ? REG_2_17 : _GEN_696; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_698 = 5'h12 == indexTagReg ? REG_2_18 : _GEN_697; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_699 = 5'h13 == indexTagReg ? REG_2_19 : _GEN_698; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_700 = 5'h14 == indexTagReg ? REG_2_20 : _GEN_699; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_701 = 5'h15 == indexTagReg ? REG_2_21 : _GEN_700; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_702 = 5'h16 == indexTagReg ? REG_2_22 : _GEN_701; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_703 = 5'h17 == indexTagReg ? REG_2_23 : _GEN_702; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_704 = 5'h18 == indexTagReg ? REG_2_24 : _GEN_703; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_705 = 5'h19 == indexTagReg ? REG_2_25 : _GEN_704; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_706 = 5'h1a == indexTagReg ? REG_2_26 : _GEN_705; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_707 = 5'h1b == indexTagReg ? REG_2_27 : _GEN_706; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_708 = 5'h1c == indexTagReg ? REG_2_28 : _GEN_707; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_709 = 5'h1d == indexTagReg ? REG_2_29 : _GEN_708; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_712 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_10_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_713 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_10_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_714 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_10_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_715 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_10_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_716 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_10_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_717 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_10_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_718 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_10_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_719 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_10_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_720 = 4'h8 == _GEN_2632 | REG_10_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_721 = 4'h9 == _GEN_2632 | REG_10_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_722 = 4'ha == _GEN_2632 | REG_10_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_723 = 4'hb == _GEN_2632 | REG_10_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_724 = 4'hc == _GEN_2632 | REG_10_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_725 = 4'hd == _GEN_2632 | REG_10_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_726 = 4'he == _GEN_2632 | REG_10_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_727 = 4'hf == _GEN_2632 | REG_10_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_728 = 5'h10 == _GEN_2648 | REG_10_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_729 = 5'h11 == _GEN_2648 | REG_10_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_730 = 5'h12 == _GEN_2648 | REG_10_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_731 = 5'h13 == _GEN_2648 | REG_10_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_732 = 5'h14 == _GEN_2648 | REG_10_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_733 = 5'h15 == _GEN_2648 | REG_10_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_734 = 5'h16 == _GEN_2648 | REG_10_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_735 = 5'h17 == _GEN_2648 | REG_10_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_736 = 5'h18 == _GEN_2648 | REG_10_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_737 = 5'h19 == _GEN_2648 | REG_10_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_738 = 5'h1a == _GEN_2648 | REG_10_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_739 = 5'h1b == _GEN_2648 | REG_10_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_740 = 5'h1c == _GEN_2648 | REG_10_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_741 = 5'h1d == _GEN_2648 | REG_10_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_742 = 5'h1e == _GEN_2648 | REG_10_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_743 = 5'h1f == _GEN_2648 | REG_10_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_744 = _GEN_2624 | REG_2_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_745 = _GEN_2625 | REG_2_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_746 = _GEN_2626 | REG_2_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_747 = _GEN_2627 | REG_2_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_748 = _GEN_2628 | REG_2_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_749 = _GEN_2629 | REG_2_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_750 = _GEN_2630 | REG_2_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_751 = _GEN_2631 | REG_2_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_752 = _GEN_2633 | REG_2_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_753 = _GEN_2635 | REG_2_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_754 = _GEN_2637 | REG_2_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_755 = _GEN_2639 | REG_2_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_756 = _GEN_2641 | REG_2_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_757 = _GEN_2643 | REG_2_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_758 = _GEN_2645 | REG_2_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_759 = _GEN_2647 | REG_2_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_760 = _GEN_2649 | REG_2_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_761 = _GEN_2651 | REG_2_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_762 = _GEN_2653 | REG_2_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_763 = _GEN_2655 | REG_2_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_764 = _GEN_2657 | REG_2_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_765 = _GEN_2659 | REG_2_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_766 = _GEN_2661 | REG_2_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_767 = _GEN_2663 | REG_2_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_768 = _GEN_2665 | REG_2_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_769 = _GEN_2667 | REG_2_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_770 = _GEN_2669 | REG_2_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_771 = _GEN_2671 | REG_2_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_772 = _GEN_2673 | REG_2_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_773 = _GEN_2675 | REG_2_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_774 = _GEN_2677 | REG_2_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_775 = _GEN_2679 | REG_2_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_776 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_777 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_778 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_779 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_780 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_781 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_782 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_783 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_2_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_784 = 4'h8 == _GEN_2632 ? 1'h0 : REG_2_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_785 = 4'h9 == _GEN_2632 ? 1'h0 : REG_2_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_786 = 4'ha == _GEN_2632 ? 1'h0 : REG_2_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_787 = 4'hb == _GEN_2632 ? 1'h0 : REG_2_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_788 = 4'hc == _GEN_2632 ? 1'h0 : REG_2_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_789 = 4'hd == _GEN_2632 ? 1'h0 : REG_2_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_790 = 4'he == _GEN_2632 ? 1'h0 : REG_2_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_791 = 4'hf == _GEN_2632 ? 1'h0 : REG_2_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_792 = 5'h10 == _GEN_2648 ? 1'h0 : REG_2_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_793 = 5'h11 == _GEN_2648 ? 1'h0 : REG_2_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_794 = 5'h12 == _GEN_2648 ? 1'h0 : REG_2_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_795 = 5'h13 == _GEN_2648 ? 1'h0 : REG_2_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_796 = 5'h14 == _GEN_2648 ? 1'h0 : REG_2_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_797 = 5'h15 == _GEN_2648 ? 1'h0 : REG_2_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_798 = 5'h16 == _GEN_2648 ? 1'h0 : REG_2_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_799 = 5'h17 == _GEN_2648 ? 1'h0 : REG_2_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_800 = 5'h18 == _GEN_2648 ? 1'h0 : REG_2_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_801 = 5'h19 == _GEN_2648 ? 1'h0 : REG_2_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_802 = 5'h1a == _GEN_2648 ? 1'h0 : REG_2_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_803 = 5'h1b == _GEN_2648 ? 1'h0 : REG_2_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_804 = 5'h1c == _GEN_2648 ? 1'h0 : REG_2_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_805 = 5'h1d == _GEN_2648 ? 1'h0 : REG_2_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_806 = 5'h1e == _GEN_2648 ? 1'h0 : REG_2_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_807 = 5'h1f == _GEN_2648 ? 1'h0 : REG_2_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_808 = updateLogic_io_cacheUpdateControl_update ? _GEN_744 : _GEN_776; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_809 = updateLogic_io_cacheUpdateControl_update ? _GEN_745 : _GEN_777; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_810 = updateLogic_io_cacheUpdateControl_update ? _GEN_746 : _GEN_778; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_811 = updateLogic_io_cacheUpdateControl_update ? _GEN_747 : _GEN_779; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_812 = updateLogic_io_cacheUpdateControl_update ? _GEN_748 : _GEN_780; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_813 = updateLogic_io_cacheUpdateControl_update ? _GEN_749 : _GEN_781; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_814 = updateLogic_io_cacheUpdateControl_update ? _GEN_750 : _GEN_782; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_815 = updateLogic_io_cacheUpdateControl_update ? _GEN_751 : _GEN_783; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_816 = updateLogic_io_cacheUpdateControl_update ? _GEN_752 : _GEN_784; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_817 = updateLogic_io_cacheUpdateControl_update ? _GEN_753 : _GEN_785; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_818 = updateLogic_io_cacheUpdateControl_update ? _GEN_754 : _GEN_786; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_819 = updateLogic_io_cacheUpdateControl_update ? _GEN_755 : _GEN_787; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_820 = updateLogic_io_cacheUpdateControl_update ? _GEN_756 : _GEN_788; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_821 = updateLogic_io_cacheUpdateControl_update ? _GEN_757 : _GEN_789; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_822 = updateLogic_io_cacheUpdateControl_update ? _GEN_758 : _GEN_790; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_823 = updateLogic_io_cacheUpdateControl_update ? _GEN_759 : _GEN_791; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_824 = updateLogic_io_cacheUpdateControl_update ? _GEN_760 : _GEN_792; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_825 = updateLogic_io_cacheUpdateControl_update ? _GEN_761 : _GEN_793; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_826 = updateLogic_io_cacheUpdateControl_update ? _GEN_762 : _GEN_794; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_827 = updateLogic_io_cacheUpdateControl_update ? _GEN_763 : _GEN_795; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_828 = updateLogic_io_cacheUpdateControl_update ? _GEN_764 : _GEN_796; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_829 = updateLogic_io_cacheUpdateControl_update ? _GEN_765 : _GEN_797; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_830 = updateLogic_io_cacheUpdateControl_update ? _GEN_766 : _GEN_798; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_831 = updateLogic_io_cacheUpdateControl_update ? _GEN_767 : _GEN_799; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_832 = updateLogic_io_cacheUpdateControl_update ? _GEN_768 : _GEN_800; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_833 = updateLogic_io_cacheUpdateControl_update ? _GEN_769 : _GEN_801; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_834 = updateLogic_io_cacheUpdateControl_update ? _GEN_770 : _GEN_802; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_835 = updateLogic_io_cacheUpdateControl_update ? _GEN_771 : _GEN_803; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_836 = updateLogic_io_cacheUpdateControl_update ? _GEN_772 : _GEN_804; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_837 = updateLogic_io_cacheUpdateControl_update ? _GEN_773 : _GEN_805; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_838 = updateLogic_io_cacheUpdateControl_update ? _GEN_774 : _GEN_806; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_839 = updateLogic_io_cacheUpdateControl_update ? _GEN_775 : _GEN_807; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_872 = _T_2 ? _GEN_808 : REG_2_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_873 = _T_2 ? _GEN_809 : REG_2_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_874 = _T_2 ? _GEN_810 : REG_2_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_875 = _T_2 ? _GEN_811 : REG_2_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_876 = _T_2 ? _GEN_812 : REG_2_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_877 = _T_2 ? _GEN_813 : REG_2_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_878 = _T_2 ? _GEN_814 : REG_2_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_879 = _T_2 ? _GEN_815 : REG_2_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_880 = _T_2 ? _GEN_816 : REG_2_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_881 = _T_2 ? _GEN_817 : REG_2_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_882 = _T_2 ? _GEN_818 : REG_2_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_883 = _T_2 ? _GEN_819 : REG_2_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_884 = _T_2 ? _GEN_820 : REG_2_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_885 = _T_2 ? _GEN_821 : REG_2_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_886 = _T_2 ? _GEN_822 : REG_2_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_887 = _T_2 ? _GEN_823 : REG_2_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_888 = _T_2 ? _GEN_824 : REG_2_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_889 = _T_2 ? _GEN_825 : REG_2_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_890 = _T_2 ? _GEN_826 : REG_2_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_891 = _T_2 ? _GEN_827 : REG_2_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_892 = _T_2 ? _GEN_828 : REG_2_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_893 = _T_2 ? _GEN_829 : REG_2_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_894 = _T_2 ? _GEN_830 : REG_2_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_895 = _T_2 ? _GEN_831 : REG_2_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_896 = _T_2 ? _GEN_832 : REG_2_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_897 = _T_2 ? _GEN_833 : REG_2_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_898 = _T_2 ? _GEN_834 : REG_2_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_899 = _T_2 ? _GEN_835 : REG_2_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_900 = _T_2 ? _GEN_836 : REG_2_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_901 = _T_2 ? _GEN_837 : REG_2_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_902 = _T_2 ? _GEN_838 : REG_2_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_903 = _T_2 ? _GEN_839 : REG_2_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_904 = _GEN_2624 | _GEN_872; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_905 = _GEN_2625 | _GEN_873; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_906 = _GEN_2626 | _GEN_874; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_907 = _GEN_2627 | _GEN_875; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_908 = _GEN_2628 | _GEN_876; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_909 = _GEN_2629 | _GEN_877; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_910 = _GEN_2630 | _GEN_878; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_911 = _GEN_2631 | _GEN_879; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_912 = _GEN_2633 | _GEN_880; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_913 = _GEN_2635 | _GEN_881; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_914 = _GEN_2637 | _GEN_882; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_915 = _GEN_2639 | _GEN_883; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_916 = _GEN_2641 | _GEN_884; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_917 = _GEN_2643 | _GEN_885; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_918 = _GEN_2645 | _GEN_886; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_919 = _GEN_2647 | _GEN_887; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_920 = _GEN_2649 | _GEN_888; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_921 = _GEN_2651 | _GEN_889; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_922 = _GEN_2653 | _GEN_890; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_923 = _GEN_2655 | _GEN_891; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_924 = _GEN_2657 | _GEN_892; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_925 = _GEN_2659 | _GEN_893; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_926 = _GEN_2661 | _GEN_894; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_927 = _GEN_2663 | _GEN_895; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_928 = _GEN_2665 | _GEN_896; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_929 = _GEN_2667 | _GEN_897; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_930 = _GEN_2669 | _GEN_898; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_931 = _GEN_2671 | _GEN_899; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_932 = _GEN_2673 | _GEN_900; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_933 = _GEN_2675 | _GEN_901; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_934 = _GEN_2677 | _GEN_902; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_935 = _GEN_2679 | _GEN_903; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_3 = MemBlock_3_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_969 = 5'h1 == indexTagReg ? REG_11_1 : REG_11_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_970 = 5'h2 == indexTagReg ? REG_11_2 : _GEN_969; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_971 = 5'h3 == indexTagReg ? REG_11_3 : _GEN_970; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_972 = 5'h4 == indexTagReg ? REG_11_4 : _GEN_971; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_973 = 5'h5 == indexTagReg ? REG_11_5 : _GEN_972; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_974 = 5'h6 == indexTagReg ? REG_11_6 : _GEN_973; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_975 = 5'h7 == indexTagReg ? REG_11_7 : _GEN_974; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_976 = 5'h8 == indexTagReg ? REG_11_8 : _GEN_975; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_977 = 5'h9 == indexTagReg ? REG_11_9 : _GEN_976; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_978 = 5'ha == indexTagReg ? REG_11_10 : _GEN_977; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_979 = 5'hb == indexTagReg ? REG_11_11 : _GEN_978; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_980 = 5'hc == indexTagReg ? REG_11_12 : _GEN_979; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_981 = 5'hd == indexTagReg ? REG_11_13 : _GEN_980; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_982 = 5'he == indexTagReg ? REG_11_14 : _GEN_981; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_983 = 5'hf == indexTagReg ? REG_11_15 : _GEN_982; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_984 = 5'h10 == indexTagReg ? REG_11_16 : _GEN_983; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_985 = 5'h11 == indexTagReg ? REG_11_17 : _GEN_984; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_986 = 5'h12 == indexTagReg ? REG_11_18 : _GEN_985; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_987 = 5'h13 == indexTagReg ? REG_11_19 : _GEN_986; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_988 = 5'h14 == indexTagReg ? REG_11_20 : _GEN_987; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_989 = 5'h15 == indexTagReg ? REG_11_21 : _GEN_988; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_990 = 5'h16 == indexTagReg ? REG_11_22 : _GEN_989; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_991 = 5'h17 == indexTagReg ? REG_11_23 : _GEN_990; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_992 = 5'h18 == indexTagReg ? REG_11_24 : _GEN_991; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_993 = 5'h19 == indexTagReg ? REG_11_25 : _GEN_992; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_994 = 5'h1a == indexTagReg ? REG_11_26 : _GEN_993; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_995 = 5'h1b == indexTagReg ? REG_11_27 : _GEN_994; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_996 = 5'h1c == indexTagReg ? REG_11_28 : _GEN_995; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_997 = 5'h1d == indexTagReg ? REG_11_29 : _GEN_996; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_998 = 5'h1e == indexTagReg ? REG_11_30 : _GEN_997; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_999 = 5'h1f == indexTagReg ? REG_11_31 : _GEN_998; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_3 = _GEN_999 & tagTagReg == readTags_3; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_1001 = 5'h1 == indexTagReg ? REG_3_1 : REG_3_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1002 = 5'h2 == indexTagReg ? REG_3_2 : _GEN_1001; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1003 = 5'h3 == indexTagReg ? REG_3_3 : _GEN_1002; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1004 = 5'h4 == indexTagReg ? REG_3_4 : _GEN_1003; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1005 = 5'h5 == indexTagReg ? REG_3_5 : _GEN_1004; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1006 = 5'h6 == indexTagReg ? REG_3_6 : _GEN_1005; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1007 = 5'h7 == indexTagReg ? REG_3_7 : _GEN_1006; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1008 = 5'h8 == indexTagReg ? REG_3_8 : _GEN_1007; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1009 = 5'h9 == indexTagReg ? REG_3_9 : _GEN_1008; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1010 = 5'ha == indexTagReg ? REG_3_10 : _GEN_1009; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1011 = 5'hb == indexTagReg ? REG_3_11 : _GEN_1010; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1012 = 5'hc == indexTagReg ? REG_3_12 : _GEN_1011; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1013 = 5'hd == indexTagReg ? REG_3_13 : _GEN_1012; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1014 = 5'he == indexTagReg ? REG_3_14 : _GEN_1013; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1015 = 5'hf == indexTagReg ? REG_3_15 : _GEN_1014; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1016 = 5'h10 == indexTagReg ? REG_3_16 : _GEN_1015; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1017 = 5'h11 == indexTagReg ? REG_3_17 : _GEN_1016; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1018 = 5'h12 == indexTagReg ? REG_3_18 : _GEN_1017; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1019 = 5'h13 == indexTagReg ? REG_3_19 : _GEN_1018; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1020 = 5'h14 == indexTagReg ? REG_3_20 : _GEN_1019; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1021 = 5'h15 == indexTagReg ? REG_3_21 : _GEN_1020; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1022 = 5'h16 == indexTagReg ? REG_3_22 : _GEN_1021; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1023 = 5'h17 == indexTagReg ? REG_3_23 : _GEN_1022; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1024 = 5'h18 == indexTagReg ? REG_3_24 : _GEN_1023; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1025 = 5'h19 == indexTagReg ? REG_3_25 : _GEN_1024; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1026 = 5'h1a == indexTagReg ? REG_3_26 : _GEN_1025; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1027 = 5'h1b == indexTagReg ? REG_3_27 : _GEN_1026; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1028 = 5'h1c == indexTagReg ? REG_3_28 : _GEN_1027; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1029 = 5'h1d == indexTagReg ? REG_3_29 : _GEN_1028; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1032 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_11_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1033 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_11_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1034 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_11_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1035 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_11_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1036 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_11_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1037 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_11_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1038 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_11_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1039 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_11_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1040 = 4'h8 == _GEN_2632 | REG_11_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1041 = 4'h9 == _GEN_2632 | REG_11_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1042 = 4'ha == _GEN_2632 | REG_11_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1043 = 4'hb == _GEN_2632 | REG_11_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1044 = 4'hc == _GEN_2632 | REG_11_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1045 = 4'hd == _GEN_2632 | REG_11_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1046 = 4'he == _GEN_2632 | REG_11_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1047 = 4'hf == _GEN_2632 | REG_11_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1048 = 5'h10 == _GEN_2648 | REG_11_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1049 = 5'h11 == _GEN_2648 | REG_11_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1050 = 5'h12 == _GEN_2648 | REG_11_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1051 = 5'h13 == _GEN_2648 | REG_11_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1052 = 5'h14 == _GEN_2648 | REG_11_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1053 = 5'h15 == _GEN_2648 | REG_11_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1054 = 5'h16 == _GEN_2648 | REG_11_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1055 = 5'h17 == _GEN_2648 | REG_11_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1056 = 5'h18 == _GEN_2648 | REG_11_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1057 = 5'h19 == _GEN_2648 | REG_11_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1058 = 5'h1a == _GEN_2648 | REG_11_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1059 = 5'h1b == _GEN_2648 | REG_11_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1060 = 5'h1c == _GEN_2648 | REG_11_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1061 = 5'h1d == _GEN_2648 | REG_11_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1062 = 5'h1e == _GEN_2648 | REG_11_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1063 = 5'h1f == _GEN_2648 | REG_11_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1064 = _GEN_2624 | REG_3_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1065 = _GEN_2625 | REG_3_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1066 = _GEN_2626 | REG_3_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1067 = _GEN_2627 | REG_3_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1068 = _GEN_2628 | REG_3_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1069 = _GEN_2629 | REG_3_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1070 = _GEN_2630 | REG_3_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1071 = _GEN_2631 | REG_3_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1072 = _GEN_2633 | REG_3_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1073 = _GEN_2635 | REG_3_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1074 = _GEN_2637 | REG_3_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1075 = _GEN_2639 | REG_3_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1076 = _GEN_2641 | REG_3_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1077 = _GEN_2643 | REG_3_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1078 = _GEN_2645 | REG_3_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1079 = _GEN_2647 | REG_3_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1080 = _GEN_2649 | REG_3_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1081 = _GEN_2651 | REG_3_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1082 = _GEN_2653 | REG_3_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1083 = _GEN_2655 | REG_3_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1084 = _GEN_2657 | REG_3_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1085 = _GEN_2659 | REG_3_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1086 = _GEN_2661 | REG_3_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1087 = _GEN_2663 | REG_3_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1088 = _GEN_2665 | REG_3_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1089 = _GEN_2667 | REG_3_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1090 = _GEN_2669 | REG_3_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1091 = _GEN_2671 | REG_3_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1092 = _GEN_2673 | REG_3_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1093 = _GEN_2675 | REG_3_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1094 = _GEN_2677 | REG_3_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1095 = _GEN_2679 | REG_3_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1096 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1097 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1098 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1099 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1100 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1101 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1102 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1103 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_3_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1104 = 4'h8 == _GEN_2632 ? 1'h0 : REG_3_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1105 = 4'h9 == _GEN_2632 ? 1'h0 : REG_3_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1106 = 4'ha == _GEN_2632 ? 1'h0 : REG_3_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1107 = 4'hb == _GEN_2632 ? 1'h0 : REG_3_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1108 = 4'hc == _GEN_2632 ? 1'h0 : REG_3_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1109 = 4'hd == _GEN_2632 ? 1'h0 : REG_3_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1110 = 4'he == _GEN_2632 ? 1'h0 : REG_3_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1111 = 4'hf == _GEN_2632 ? 1'h0 : REG_3_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1112 = 5'h10 == _GEN_2648 ? 1'h0 : REG_3_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1113 = 5'h11 == _GEN_2648 ? 1'h0 : REG_3_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1114 = 5'h12 == _GEN_2648 ? 1'h0 : REG_3_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1115 = 5'h13 == _GEN_2648 ? 1'h0 : REG_3_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1116 = 5'h14 == _GEN_2648 ? 1'h0 : REG_3_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1117 = 5'h15 == _GEN_2648 ? 1'h0 : REG_3_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1118 = 5'h16 == _GEN_2648 ? 1'h0 : REG_3_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1119 = 5'h17 == _GEN_2648 ? 1'h0 : REG_3_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1120 = 5'h18 == _GEN_2648 ? 1'h0 : REG_3_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1121 = 5'h19 == _GEN_2648 ? 1'h0 : REG_3_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1122 = 5'h1a == _GEN_2648 ? 1'h0 : REG_3_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1123 = 5'h1b == _GEN_2648 ? 1'h0 : REG_3_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1124 = 5'h1c == _GEN_2648 ? 1'h0 : REG_3_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1125 = 5'h1d == _GEN_2648 ? 1'h0 : REG_3_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1126 = 5'h1e == _GEN_2648 ? 1'h0 : REG_3_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1127 = 5'h1f == _GEN_2648 ? 1'h0 : REG_3_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1128 = updateLogic_io_cacheUpdateControl_update ? _GEN_1064 : _GEN_1096; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1129 = updateLogic_io_cacheUpdateControl_update ? _GEN_1065 : _GEN_1097; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1130 = updateLogic_io_cacheUpdateControl_update ? _GEN_1066 : _GEN_1098; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1131 = updateLogic_io_cacheUpdateControl_update ? _GEN_1067 : _GEN_1099; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1132 = updateLogic_io_cacheUpdateControl_update ? _GEN_1068 : _GEN_1100; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1133 = updateLogic_io_cacheUpdateControl_update ? _GEN_1069 : _GEN_1101; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1134 = updateLogic_io_cacheUpdateControl_update ? _GEN_1070 : _GEN_1102; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1135 = updateLogic_io_cacheUpdateControl_update ? _GEN_1071 : _GEN_1103; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1136 = updateLogic_io_cacheUpdateControl_update ? _GEN_1072 : _GEN_1104; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1137 = updateLogic_io_cacheUpdateControl_update ? _GEN_1073 : _GEN_1105; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1138 = updateLogic_io_cacheUpdateControl_update ? _GEN_1074 : _GEN_1106; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1139 = updateLogic_io_cacheUpdateControl_update ? _GEN_1075 : _GEN_1107; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1140 = updateLogic_io_cacheUpdateControl_update ? _GEN_1076 : _GEN_1108; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1141 = updateLogic_io_cacheUpdateControl_update ? _GEN_1077 : _GEN_1109; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1142 = updateLogic_io_cacheUpdateControl_update ? _GEN_1078 : _GEN_1110; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1143 = updateLogic_io_cacheUpdateControl_update ? _GEN_1079 : _GEN_1111; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1144 = updateLogic_io_cacheUpdateControl_update ? _GEN_1080 : _GEN_1112; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1145 = updateLogic_io_cacheUpdateControl_update ? _GEN_1081 : _GEN_1113; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1146 = updateLogic_io_cacheUpdateControl_update ? _GEN_1082 : _GEN_1114; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1147 = updateLogic_io_cacheUpdateControl_update ? _GEN_1083 : _GEN_1115; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1148 = updateLogic_io_cacheUpdateControl_update ? _GEN_1084 : _GEN_1116; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1149 = updateLogic_io_cacheUpdateControl_update ? _GEN_1085 : _GEN_1117; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1150 = updateLogic_io_cacheUpdateControl_update ? _GEN_1086 : _GEN_1118; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1151 = updateLogic_io_cacheUpdateControl_update ? _GEN_1087 : _GEN_1119; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1152 = updateLogic_io_cacheUpdateControl_update ? _GEN_1088 : _GEN_1120; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1153 = updateLogic_io_cacheUpdateControl_update ? _GEN_1089 : _GEN_1121; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1154 = updateLogic_io_cacheUpdateControl_update ? _GEN_1090 : _GEN_1122; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1155 = updateLogic_io_cacheUpdateControl_update ? _GEN_1091 : _GEN_1123; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1156 = updateLogic_io_cacheUpdateControl_update ? _GEN_1092 : _GEN_1124; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1157 = updateLogic_io_cacheUpdateControl_update ? _GEN_1093 : _GEN_1125; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1158 = updateLogic_io_cacheUpdateControl_update ? _GEN_1094 : _GEN_1126; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1159 = updateLogic_io_cacheUpdateControl_update ? _GEN_1095 : _GEN_1127; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1192 = _T_3 ? _GEN_1128 : REG_3_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1193 = _T_3 ? _GEN_1129 : REG_3_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1194 = _T_3 ? _GEN_1130 : REG_3_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1195 = _T_3 ? _GEN_1131 : REG_3_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1196 = _T_3 ? _GEN_1132 : REG_3_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1197 = _T_3 ? _GEN_1133 : REG_3_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1198 = _T_3 ? _GEN_1134 : REG_3_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1199 = _T_3 ? _GEN_1135 : REG_3_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1200 = _T_3 ? _GEN_1136 : REG_3_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1201 = _T_3 ? _GEN_1137 : REG_3_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1202 = _T_3 ? _GEN_1138 : REG_3_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1203 = _T_3 ? _GEN_1139 : REG_3_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1204 = _T_3 ? _GEN_1140 : REG_3_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1205 = _T_3 ? _GEN_1141 : REG_3_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1206 = _T_3 ? _GEN_1142 : REG_3_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1207 = _T_3 ? _GEN_1143 : REG_3_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1208 = _T_3 ? _GEN_1144 : REG_3_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1209 = _T_3 ? _GEN_1145 : REG_3_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1210 = _T_3 ? _GEN_1146 : REG_3_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1211 = _T_3 ? _GEN_1147 : REG_3_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1212 = _T_3 ? _GEN_1148 : REG_3_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1213 = _T_3 ? _GEN_1149 : REG_3_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1214 = _T_3 ? _GEN_1150 : REG_3_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1215 = _T_3 ? _GEN_1151 : REG_3_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1216 = _T_3 ? _GEN_1152 : REG_3_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1217 = _T_3 ? _GEN_1153 : REG_3_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1218 = _T_3 ? _GEN_1154 : REG_3_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1219 = _T_3 ? _GEN_1155 : REG_3_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1220 = _T_3 ? _GEN_1156 : REG_3_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1221 = _T_3 ? _GEN_1157 : REG_3_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1222 = _T_3 ? _GEN_1158 : REG_3_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1223 = _T_3 ? _GEN_1159 : REG_3_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1224 = _GEN_2624 | _GEN_1192; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1225 = _GEN_2625 | _GEN_1193; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1226 = _GEN_2626 | _GEN_1194; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1227 = _GEN_2627 | _GEN_1195; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1228 = _GEN_2628 | _GEN_1196; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1229 = _GEN_2629 | _GEN_1197; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1230 = _GEN_2630 | _GEN_1198; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1231 = _GEN_2631 | _GEN_1199; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1232 = _GEN_2633 | _GEN_1200; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1233 = _GEN_2635 | _GEN_1201; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1234 = _GEN_2637 | _GEN_1202; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1235 = _GEN_2639 | _GEN_1203; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1236 = _GEN_2641 | _GEN_1204; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1237 = _GEN_2643 | _GEN_1205; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1238 = _GEN_2645 | _GEN_1206; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1239 = _GEN_2647 | _GEN_1207; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1240 = _GEN_2649 | _GEN_1208; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1241 = _GEN_2651 | _GEN_1209; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1242 = _GEN_2653 | _GEN_1210; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1243 = _GEN_2655 | _GEN_1211; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1244 = _GEN_2657 | _GEN_1212; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1245 = _GEN_2659 | _GEN_1213; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1246 = _GEN_2661 | _GEN_1214; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1247 = _GEN_2663 | _GEN_1215; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1248 = _GEN_2665 | _GEN_1216; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1249 = _GEN_2667 | _GEN_1217; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1250 = _GEN_2669 | _GEN_1218; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1251 = _GEN_2671 | _GEN_1219; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1252 = _GEN_2673 | _GEN_1220; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1253 = _GEN_2675 | _GEN_1221; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1254 = _GEN_2677 | _GEN_1222; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1255 = _GEN_2679 | _GEN_1223; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_4 = MemBlock_4_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_1289 = 5'h1 == indexTagReg ? REG_12_1 : REG_12_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1290 = 5'h2 == indexTagReg ? REG_12_2 : _GEN_1289; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1291 = 5'h3 == indexTagReg ? REG_12_3 : _GEN_1290; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1292 = 5'h4 == indexTagReg ? REG_12_4 : _GEN_1291; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1293 = 5'h5 == indexTagReg ? REG_12_5 : _GEN_1292; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1294 = 5'h6 == indexTagReg ? REG_12_6 : _GEN_1293; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1295 = 5'h7 == indexTagReg ? REG_12_7 : _GEN_1294; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1296 = 5'h8 == indexTagReg ? REG_12_8 : _GEN_1295; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1297 = 5'h9 == indexTagReg ? REG_12_9 : _GEN_1296; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1298 = 5'ha == indexTagReg ? REG_12_10 : _GEN_1297; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1299 = 5'hb == indexTagReg ? REG_12_11 : _GEN_1298; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1300 = 5'hc == indexTagReg ? REG_12_12 : _GEN_1299; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1301 = 5'hd == indexTagReg ? REG_12_13 : _GEN_1300; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1302 = 5'he == indexTagReg ? REG_12_14 : _GEN_1301; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1303 = 5'hf == indexTagReg ? REG_12_15 : _GEN_1302; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1304 = 5'h10 == indexTagReg ? REG_12_16 : _GEN_1303; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1305 = 5'h11 == indexTagReg ? REG_12_17 : _GEN_1304; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1306 = 5'h12 == indexTagReg ? REG_12_18 : _GEN_1305; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1307 = 5'h13 == indexTagReg ? REG_12_19 : _GEN_1306; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1308 = 5'h14 == indexTagReg ? REG_12_20 : _GEN_1307; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1309 = 5'h15 == indexTagReg ? REG_12_21 : _GEN_1308; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1310 = 5'h16 == indexTagReg ? REG_12_22 : _GEN_1309; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1311 = 5'h17 == indexTagReg ? REG_12_23 : _GEN_1310; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1312 = 5'h18 == indexTagReg ? REG_12_24 : _GEN_1311; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1313 = 5'h19 == indexTagReg ? REG_12_25 : _GEN_1312; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1314 = 5'h1a == indexTagReg ? REG_12_26 : _GEN_1313; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1315 = 5'h1b == indexTagReg ? REG_12_27 : _GEN_1314; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1316 = 5'h1c == indexTagReg ? REG_12_28 : _GEN_1315; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1317 = 5'h1d == indexTagReg ? REG_12_29 : _GEN_1316; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1318 = 5'h1e == indexTagReg ? REG_12_30 : _GEN_1317; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1319 = 5'h1f == indexTagReg ? REG_12_31 : _GEN_1318; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_4 = _GEN_1319 & tagTagReg == readTags_4; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_1321 = 5'h1 == indexTagReg ? REG_4_1 : REG_4_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1322 = 5'h2 == indexTagReg ? REG_4_2 : _GEN_1321; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1323 = 5'h3 == indexTagReg ? REG_4_3 : _GEN_1322; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1324 = 5'h4 == indexTagReg ? REG_4_4 : _GEN_1323; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1325 = 5'h5 == indexTagReg ? REG_4_5 : _GEN_1324; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1326 = 5'h6 == indexTagReg ? REG_4_6 : _GEN_1325; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1327 = 5'h7 == indexTagReg ? REG_4_7 : _GEN_1326; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1328 = 5'h8 == indexTagReg ? REG_4_8 : _GEN_1327; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1329 = 5'h9 == indexTagReg ? REG_4_9 : _GEN_1328; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1330 = 5'ha == indexTagReg ? REG_4_10 : _GEN_1329; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1331 = 5'hb == indexTagReg ? REG_4_11 : _GEN_1330; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1332 = 5'hc == indexTagReg ? REG_4_12 : _GEN_1331; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1333 = 5'hd == indexTagReg ? REG_4_13 : _GEN_1332; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1334 = 5'he == indexTagReg ? REG_4_14 : _GEN_1333; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1335 = 5'hf == indexTagReg ? REG_4_15 : _GEN_1334; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1336 = 5'h10 == indexTagReg ? REG_4_16 : _GEN_1335; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1337 = 5'h11 == indexTagReg ? REG_4_17 : _GEN_1336; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1338 = 5'h12 == indexTagReg ? REG_4_18 : _GEN_1337; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1339 = 5'h13 == indexTagReg ? REG_4_19 : _GEN_1338; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1340 = 5'h14 == indexTagReg ? REG_4_20 : _GEN_1339; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1341 = 5'h15 == indexTagReg ? REG_4_21 : _GEN_1340; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1342 = 5'h16 == indexTagReg ? REG_4_22 : _GEN_1341; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1343 = 5'h17 == indexTagReg ? REG_4_23 : _GEN_1342; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1344 = 5'h18 == indexTagReg ? REG_4_24 : _GEN_1343; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1345 = 5'h19 == indexTagReg ? REG_4_25 : _GEN_1344; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1346 = 5'h1a == indexTagReg ? REG_4_26 : _GEN_1345; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1347 = 5'h1b == indexTagReg ? REG_4_27 : _GEN_1346; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1348 = 5'h1c == indexTagReg ? REG_4_28 : _GEN_1347; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1349 = 5'h1d == indexTagReg ? REG_4_29 : _GEN_1348; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1352 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_12_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1353 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_12_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1354 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_12_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1355 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_12_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1356 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_12_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1357 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_12_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1358 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_12_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1359 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_12_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1360 = 4'h8 == _GEN_2632 | REG_12_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1361 = 4'h9 == _GEN_2632 | REG_12_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1362 = 4'ha == _GEN_2632 | REG_12_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1363 = 4'hb == _GEN_2632 | REG_12_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1364 = 4'hc == _GEN_2632 | REG_12_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1365 = 4'hd == _GEN_2632 | REG_12_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1366 = 4'he == _GEN_2632 | REG_12_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1367 = 4'hf == _GEN_2632 | REG_12_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1368 = 5'h10 == _GEN_2648 | REG_12_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1369 = 5'h11 == _GEN_2648 | REG_12_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1370 = 5'h12 == _GEN_2648 | REG_12_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1371 = 5'h13 == _GEN_2648 | REG_12_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1372 = 5'h14 == _GEN_2648 | REG_12_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1373 = 5'h15 == _GEN_2648 | REG_12_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1374 = 5'h16 == _GEN_2648 | REG_12_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1375 = 5'h17 == _GEN_2648 | REG_12_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1376 = 5'h18 == _GEN_2648 | REG_12_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1377 = 5'h19 == _GEN_2648 | REG_12_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1378 = 5'h1a == _GEN_2648 | REG_12_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1379 = 5'h1b == _GEN_2648 | REG_12_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1380 = 5'h1c == _GEN_2648 | REG_12_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1381 = 5'h1d == _GEN_2648 | REG_12_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1382 = 5'h1e == _GEN_2648 | REG_12_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1383 = 5'h1f == _GEN_2648 | REG_12_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1384 = _GEN_2624 | REG_4_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1385 = _GEN_2625 | REG_4_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1386 = _GEN_2626 | REG_4_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1387 = _GEN_2627 | REG_4_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1388 = _GEN_2628 | REG_4_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1389 = _GEN_2629 | REG_4_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1390 = _GEN_2630 | REG_4_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1391 = _GEN_2631 | REG_4_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1392 = _GEN_2633 | REG_4_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1393 = _GEN_2635 | REG_4_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1394 = _GEN_2637 | REG_4_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1395 = _GEN_2639 | REG_4_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1396 = _GEN_2641 | REG_4_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1397 = _GEN_2643 | REG_4_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1398 = _GEN_2645 | REG_4_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1399 = _GEN_2647 | REG_4_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1400 = _GEN_2649 | REG_4_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1401 = _GEN_2651 | REG_4_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1402 = _GEN_2653 | REG_4_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1403 = _GEN_2655 | REG_4_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1404 = _GEN_2657 | REG_4_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1405 = _GEN_2659 | REG_4_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1406 = _GEN_2661 | REG_4_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1407 = _GEN_2663 | REG_4_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1408 = _GEN_2665 | REG_4_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1409 = _GEN_2667 | REG_4_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1410 = _GEN_2669 | REG_4_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1411 = _GEN_2671 | REG_4_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1412 = _GEN_2673 | REG_4_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1413 = _GEN_2675 | REG_4_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1414 = _GEN_2677 | REG_4_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1415 = _GEN_2679 | REG_4_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1416 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1417 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1418 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1419 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1420 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1421 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1422 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1423 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_4_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1424 = 4'h8 == _GEN_2632 ? 1'h0 : REG_4_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1425 = 4'h9 == _GEN_2632 ? 1'h0 : REG_4_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1426 = 4'ha == _GEN_2632 ? 1'h0 : REG_4_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1427 = 4'hb == _GEN_2632 ? 1'h0 : REG_4_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1428 = 4'hc == _GEN_2632 ? 1'h0 : REG_4_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1429 = 4'hd == _GEN_2632 ? 1'h0 : REG_4_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1430 = 4'he == _GEN_2632 ? 1'h0 : REG_4_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1431 = 4'hf == _GEN_2632 ? 1'h0 : REG_4_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1432 = 5'h10 == _GEN_2648 ? 1'h0 : REG_4_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1433 = 5'h11 == _GEN_2648 ? 1'h0 : REG_4_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1434 = 5'h12 == _GEN_2648 ? 1'h0 : REG_4_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1435 = 5'h13 == _GEN_2648 ? 1'h0 : REG_4_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1436 = 5'h14 == _GEN_2648 ? 1'h0 : REG_4_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1437 = 5'h15 == _GEN_2648 ? 1'h0 : REG_4_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1438 = 5'h16 == _GEN_2648 ? 1'h0 : REG_4_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1439 = 5'h17 == _GEN_2648 ? 1'h0 : REG_4_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1440 = 5'h18 == _GEN_2648 ? 1'h0 : REG_4_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1441 = 5'h19 == _GEN_2648 ? 1'h0 : REG_4_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1442 = 5'h1a == _GEN_2648 ? 1'h0 : REG_4_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1443 = 5'h1b == _GEN_2648 ? 1'h0 : REG_4_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1444 = 5'h1c == _GEN_2648 ? 1'h0 : REG_4_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1445 = 5'h1d == _GEN_2648 ? 1'h0 : REG_4_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1446 = 5'h1e == _GEN_2648 ? 1'h0 : REG_4_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1447 = 5'h1f == _GEN_2648 ? 1'h0 : REG_4_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1448 = updateLogic_io_cacheUpdateControl_update ? _GEN_1384 : _GEN_1416; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1449 = updateLogic_io_cacheUpdateControl_update ? _GEN_1385 : _GEN_1417; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1450 = updateLogic_io_cacheUpdateControl_update ? _GEN_1386 : _GEN_1418; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1451 = updateLogic_io_cacheUpdateControl_update ? _GEN_1387 : _GEN_1419; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1452 = updateLogic_io_cacheUpdateControl_update ? _GEN_1388 : _GEN_1420; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1453 = updateLogic_io_cacheUpdateControl_update ? _GEN_1389 : _GEN_1421; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1454 = updateLogic_io_cacheUpdateControl_update ? _GEN_1390 : _GEN_1422; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1455 = updateLogic_io_cacheUpdateControl_update ? _GEN_1391 : _GEN_1423; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1456 = updateLogic_io_cacheUpdateControl_update ? _GEN_1392 : _GEN_1424; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1457 = updateLogic_io_cacheUpdateControl_update ? _GEN_1393 : _GEN_1425; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1458 = updateLogic_io_cacheUpdateControl_update ? _GEN_1394 : _GEN_1426; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1459 = updateLogic_io_cacheUpdateControl_update ? _GEN_1395 : _GEN_1427; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1460 = updateLogic_io_cacheUpdateControl_update ? _GEN_1396 : _GEN_1428; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1461 = updateLogic_io_cacheUpdateControl_update ? _GEN_1397 : _GEN_1429; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1462 = updateLogic_io_cacheUpdateControl_update ? _GEN_1398 : _GEN_1430; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1463 = updateLogic_io_cacheUpdateControl_update ? _GEN_1399 : _GEN_1431; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1464 = updateLogic_io_cacheUpdateControl_update ? _GEN_1400 : _GEN_1432; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1465 = updateLogic_io_cacheUpdateControl_update ? _GEN_1401 : _GEN_1433; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1466 = updateLogic_io_cacheUpdateControl_update ? _GEN_1402 : _GEN_1434; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1467 = updateLogic_io_cacheUpdateControl_update ? _GEN_1403 : _GEN_1435; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1468 = updateLogic_io_cacheUpdateControl_update ? _GEN_1404 : _GEN_1436; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1469 = updateLogic_io_cacheUpdateControl_update ? _GEN_1405 : _GEN_1437; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1470 = updateLogic_io_cacheUpdateControl_update ? _GEN_1406 : _GEN_1438; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1471 = updateLogic_io_cacheUpdateControl_update ? _GEN_1407 : _GEN_1439; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1472 = updateLogic_io_cacheUpdateControl_update ? _GEN_1408 : _GEN_1440; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1473 = updateLogic_io_cacheUpdateControl_update ? _GEN_1409 : _GEN_1441; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1474 = updateLogic_io_cacheUpdateControl_update ? _GEN_1410 : _GEN_1442; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1475 = updateLogic_io_cacheUpdateControl_update ? _GEN_1411 : _GEN_1443; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1476 = updateLogic_io_cacheUpdateControl_update ? _GEN_1412 : _GEN_1444; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1477 = updateLogic_io_cacheUpdateControl_update ? _GEN_1413 : _GEN_1445; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1478 = updateLogic_io_cacheUpdateControl_update ? _GEN_1414 : _GEN_1446; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1479 = updateLogic_io_cacheUpdateControl_update ? _GEN_1415 : _GEN_1447; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1512 = _T_4 ? _GEN_1448 : REG_4_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1513 = _T_4 ? _GEN_1449 : REG_4_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1514 = _T_4 ? _GEN_1450 : REG_4_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1515 = _T_4 ? _GEN_1451 : REG_4_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1516 = _T_4 ? _GEN_1452 : REG_4_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1517 = _T_4 ? _GEN_1453 : REG_4_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1518 = _T_4 ? _GEN_1454 : REG_4_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1519 = _T_4 ? _GEN_1455 : REG_4_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1520 = _T_4 ? _GEN_1456 : REG_4_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1521 = _T_4 ? _GEN_1457 : REG_4_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1522 = _T_4 ? _GEN_1458 : REG_4_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1523 = _T_4 ? _GEN_1459 : REG_4_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1524 = _T_4 ? _GEN_1460 : REG_4_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1525 = _T_4 ? _GEN_1461 : REG_4_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1526 = _T_4 ? _GEN_1462 : REG_4_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1527 = _T_4 ? _GEN_1463 : REG_4_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1528 = _T_4 ? _GEN_1464 : REG_4_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1529 = _T_4 ? _GEN_1465 : REG_4_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1530 = _T_4 ? _GEN_1466 : REG_4_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1531 = _T_4 ? _GEN_1467 : REG_4_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1532 = _T_4 ? _GEN_1468 : REG_4_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1533 = _T_4 ? _GEN_1469 : REG_4_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1534 = _T_4 ? _GEN_1470 : REG_4_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1535 = _T_4 ? _GEN_1471 : REG_4_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1536 = _T_4 ? _GEN_1472 : REG_4_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1537 = _T_4 ? _GEN_1473 : REG_4_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1538 = _T_4 ? _GEN_1474 : REG_4_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1539 = _T_4 ? _GEN_1475 : REG_4_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1540 = _T_4 ? _GEN_1476 : REG_4_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1541 = _T_4 ? _GEN_1477 : REG_4_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1542 = _T_4 ? _GEN_1478 : REG_4_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1543 = _T_4 ? _GEN_1479 : REG_4_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1544 = _GEN_2624 | _GEN_1512; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1545 = _GEN_2625 | _GEN_1513; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1546 = _GEN_2626 | _GEN_1514; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1547 = _GEN_2627 | _GEN_1515; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1548 = _GEN_2628 | _GEN_1516; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1549 = _GEN_2629 | _GEN_1517; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1550 = _GEN_2630 | _GEN_1518; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1551 = _GEN_2631 | _GEN_1519; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1552 = _GEN_2633 | _GEN_1520; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1553 = _GEN_2635 | _GEN_1521; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1554 = _GEN_2637 | _GEN_1522; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1555 = _GEN_2639 | _GEN_1523; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1556 = _GEN_2641 | _GEN_1524; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1557 = _GEN_2643 | _GEN_1525; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1558 = _GEN_2645 | _GEN_1526; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1559 = _GEN_2647 | _GEN_1527; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1560 = _GEN_2649 | _GEN_1528; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1561 = _GEN_2651 | _GEN_1529; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1562 = _GEN_2653 | _GEN_1530; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1563 = _GEN_2655 | _GEN_1531; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1564 = _GEN_2657 | _GEN_1532; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1565 = _GEN_2659 | _GEN_1533; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1566 = _GEN_2661 | _GEN_1534; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1567 = _GEN_2663 | _GEN_1535; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1568 = _GEN_2665 | _GEN_1536; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1569 = _GEN_2667 | _GEN_1537; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1570 = _GEN_2669 | _GEN_1538; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1571 = _GEN_2671 | _GEN_1539; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1572 = _GEN_2673 | _GEN_1540; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1573 = _GEN_2675 | _GEN_1541; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1574 = _GEN_2677 | _GEN_1542; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1575 = _GEN_2679 | _GEN_1543; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_5 = MemBlock_5_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_1609 = 5'h1 == indexTagReg ? REG_13_1 : REG_13_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1610 = 5'h2 == indexTagReg ? REG_13_2 : _GEN_1609; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1611 = 5'h3 == indexTagReg ? REG_13_3 : _GEN_1610; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1612 = 5'h4 == indexTagReg ? REG_13_4 : _GEN_1611; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1613 = 5'h5 == indexTagReg ? REG_13_5 : _GEN_1612; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1614 = 5'h6 == indexTagReg ? REG_13_6 : _GEN_1613; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1615 = 5'h7 == indexTagReg ? REG_13_7 : _GEN_1614; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1616 = 5'h8 == indexTagReg ? REG_13_8 : _GEN_1615; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1617 = 5'h9 == indexTagReg ? REG_13_9 : _GEN_1616; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1618 = 5'ha == indexTagReg ? REG_13_10 : _GEN_1617; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1619 = 5'hb == indexTagReg ? REG_13_11 : _GEN_1618; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1620 = 5'hc == indexTagReg ? REG_13_12 : _GEN_1619; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1621 = 5'hd == indexTagReg ? REG_13_13 : _GEN_1620; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1622 = 5'he == indexTagReg ? REG_13_14 : _GEN_1621; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1623 = 5'hf == indexTagReg ? REG_13_15 : _GEN_1622; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1624 = 5'h10 == indexTagReg ? REG_13_16 : _GEN_1623; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1625 = 5'h11 == indexTagReg ? REG_13_17 : _GEN_1624; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1626 = 5'h12 == indexTagReg ? REG_13_18 : _GEN_1625; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1627 = 5'h13 == indexTagReg ? REG_13_19 : _GEN_1626; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1628 = 5'h14 == indexTagReg ? REG_13_20 : _GEN_1627; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1629 = 5'h15 == indexTagReg ? REG_13_21 : _GEN_1628; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1630 = 5'h16 == indexTagReg ? REG_13_22 : _GEN_1629; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1631 = 5'h17 == indexTagReg ? REG_13_23 : _GEN_1630; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1632 = 5'h18 == indexTagReg ? REG_13_24 : _GEN_1631; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1633 = 5'h19 == indexTagReg ? REG_13_25 : _GEN_1632; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1634 = 5'h1a == indexTagReg ? REG_13_26 : _GEN_1633; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1635 = 5'h1b == indexTagReg ? REG_13_27 : _GEN_1634; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1636 = 5'h1c == indexTagReg ? REG_13_28 : _GEN_1635; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1637 = 5'h1d == indexTagReg ? REG_13_29 : _GEN_1636; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1638 = 5'h1e == indexTagReg ? REG_13_30 : _GEN_1637; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1639 = 5'h1f == indexTagReg ? REG_13_31 : _GEN_1638; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_5 = _GEN_1639 & tagTagReg == readTags_5; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_1641 = 5'h1 == indexTagReg ? REG_5_1 : REG_5_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1642 = 5'h2 == indexTagReg ? REG_5_2 : _GEN_1641; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1643 = 5'h3 == indexTagReg ? REG_5_3 : _GEN_1642; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1644 = 5'h4 == indexTagReg ? REG_5_4 : _GEN_1643; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1645 = 5'h5 == indexTagReg ? REG_5_5 : _GEN_1644; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1646 = 5'h6 == indexTagReg ? REG_5_6 : _GEN_1645; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1647 = 5'h7 == indexTagReg ? REG_5_7 : _GEN_1646; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1648 = 5'h8 == indexTagReg ? REG_5_8 : _GEN_1647; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1649 = 5'h9 == indexTagReg ? REG_5_9 : _GEN_1648; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1650 = 5'ha == indexTagReg ? REG_5_10 : _GEN_1649; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1651 = 5'hb == indexTagReg ? REG_5_11 : _GEN_1650; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1652 = 5'hc == indexTagReg ? REG_5_12 : _GEN_1651; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1653 = 5'hd == indexTagReg ? REG_5_13 : _GEN_1652; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1654 = 5'he == indexTagReg ? REG_5_14 : _GEN_1653; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1655 = 5'hf == indexTagReg ? REG_5_15 : _GEN_1654; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1656 = 5'h10 == indexTagReg ? REG_5_16 : _GEN_1655; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1657 = 5'h11 == indexTagReg ? REG_5_17 : _GEN_1656; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1658 = 5'h12 == indexTagReg ? REG_5_18 : _GEN_1657; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1659 = 5'h13 == indexTagReg ? REG_5_19 : _GEN_1658; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1660 = 5'h14 == indexTagReg ? REG_5_20 : _GEN_1659; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1661 = 5'h15 == indexTagReg ? REG_5_21 : _GEN_1660; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1662 = 5'h16 == indexTagReg ? REG_5_22 : _GEN_1661; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1663 = 5'h17 == indexTagReg ? REG_5_23 : _GEN_1662; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1664 = 5'h18 == indexTagReg ? REG_5_24 : _GEN_1663; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1665 = 5'h19 == indexTagReg ? REG_5_25 : _GEN_1664; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1666 = 5'h1a == indexTagReg ? REG_5_26 : _GEN_1665; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1667 = 5'h1b == indexTagReg ? REG_5_27 : _GEN_1666; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1668 = 5'h1c == indexTagReg ? REG_5_28 : _GEN_1667; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1669 = 5'h1d == indexTagReg ? REG_5_29 : _GEN_1668; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1672 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_13_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1673 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_13_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1674 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_13_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1675 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_13_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1676 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_13_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1677 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_13_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1678 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_13_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1679 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_13_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1680 = 4'h8 == _GEN_2632 | REG_13_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1681 = 4'h9 == _GEN_2632 | REG_13_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1682 = 4'ha == _GEN_2632 | REG_13_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1683 = 4'hb == _GEN_2632 | REG_13_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1684 = 4'hc == _GEN_2632 | REG_13_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1685 = 4'hd == _GEN_2632 | REG_13_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1686 = 4'he == _GEN_2632 | REG_13_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1687 = 4'hf == _GEN_2632 | REG_13_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1688 = 5'h10 == _GEN_2648 | REG_13_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1689 = 5'h11 == _GEN_2648 | REG_13_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1690 = 5'h12 == _GEN_2648 | REG_13_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1691 = 5'h13 == _GEN_2648 | REG_13_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1692 = 5'h14 == _GEN_2648 | REG_13_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1693 = 5'h15 == _GEN_2648 | REG_13_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1694 = 5'h16 == _GEN_2648 | REG_13_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1695 = 5'h17 == _GEN_2648 | REG_13_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1696 = 5'h18 == _GEN_2648 | REG_13_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1697 = 5'h19 == _GEN_2648 | REG_13_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1698 = 5'h1a == _GEN_2648 | REG_13_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1699 = 5'h1b == _GEN_2648 | REG_13_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1700 = 5'h1c == _GEN_2648 | REG_13_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1701 = 5'h1d == _GEN_2648 | REG_13_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1702 = 5'h1e == _GEN_2648 | REG_13_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1703 = 5'h1f == _GEN_2648 | REG_13_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1704 = _GEN_2624 | REG_5_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1705 = _GEN_2625 | REG_5_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1706 = _GEN_2626 | REG_5_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1707 = _GEN_2627 | REG_5_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1708 = _GEN_2628 | REG_5_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1709 = _GEN_2629 | REG_5_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1710 = _GEN_2630 | REG_5_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1711 = _GEN_2631 | REG_5_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1712 = _GEN_2633 | REG_5_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1713 = _GEN_2635 | REG_5_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1714 = _GEN_2637 | REG_5_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1715 = _GEN_2639 | REG_5_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1716 = _GEN_2641 | REG_5_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1717 = _GEN_2643 | REG_5_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1718 = _GEN_2645 | REG_5_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1719 = _GEN_2647 | REG_5_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1720 = _GEN_2649 | REG_5_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1721 = _GEN_2651 | REG_5_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1722 = _GEN_2653 | REG_5_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1723 = _GEN_2655 | REG_5_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1724 = _GEN_2657 | REG_5_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1725 = _GEN_2659 | REG_5_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1726 = _GEN_2661 | REG_5_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1727 = _GEN_2663 | REG_5_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1728 = _GEN_2665 | REG_5_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1729 = _GEN_2667 | REG_5_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1730 = _GEN_2669 | REG_5_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1731 = _GEN_2671 | REG_5_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1732 = _GEN_2673 | REG_5_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1733 = _GEN_2675 | REG_5_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1734 = _GEN_2677 | REG_5_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1735 = _GEN_2679 | REG_5_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_1736 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1737 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1738 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1739 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1740 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1741 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1742 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1743 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_5_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1744 = 4'h8 == _GEN_2632 ? 1'h0 : REG_5_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1745 = 4'h9 == _GEN_2632 ? 1'h0 : REG_5_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1746 = 4'ha == _GEN_2632 ? 1'h0 : REG_5_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1747 = 4'hb == _GEN_2632 ? 1'h0 : REG_5_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1748 = 4'hc == _GEN_2632 ? 1'h0 : REG_5_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1749 = 4'hd == _GEN_2632 ? 1'h0 : REG_5_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1750 = 4'he == _GEN_2632 ? 1'h0 : REG_5_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1751 = 4'hf == _GEN_2632 ? 1'h0 : REG_5_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1752 = 5'h10 == _GEN_2648 ? 1'h0 : REG_5_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1753 = 5'h11 == _GEN_2648 ? 1'h0 : REG_5_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1754 = 5'h12 == _GEN_2648 ? 1'h0 : REG_5_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1755 = 5'h13 == _GEN_2648 ? 1'h0 : REG_5_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1756 = 5'h14 == _GEN_2648 ? 1'h0 : REG_5_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1757 = 5'h15 == _GEN_2648 ? 1'h0 : REG_5_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1758 = 5'h16 == _GEN_2648 ? 1'h0 : REG_5_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1759 = 5'h17 == _GEN_2648 ? 1'h0 : REG_5_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1760 = 5'h18 == _GEN_2648 ? 1'h0 : REG_5_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1761 = 5'h19 == _GEN_2648 ? 1'h0 : REG_5_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1762 = 5'h1a == _GEN_2648 ? 1'h0 : REG_5_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1763 = 5'h1b == _GEN_2648 ? 1'h0 : REG_5_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1764 = 5'h1c == _GEN_2648 ? 1'h0 : REG_5_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1765 = 5'h1d == _GEN_2648 ? 1'h0 : REG_5_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1766 = 5'h1e == _GEN_2648 ? 1'h0 : REG_5_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1767 = 5'h1f == _GEN_2648 ? 1'h0 : REG_5_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_1768 = updateLogic_io_cacheUpdateControl_update ? _GEN_1704 : _GEN_1736; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1769 = updateLogic_io_cacheUpdateControl_update ? _GEN_1705 : _GEN_1737; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1770 = updateLogic_io_cacheUpdateControl_update ? _GEN_1706 : _GEN_1738; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1771 = updateLogic_io_cacheUpdateControl_update ? _GEN_1707 : _GEN_1739; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1772 = updateLogic_io_cacheUpdateControl_update ? _GEN_1708 : _GEN_1740; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1773 = updateLogic_io_cacheUpdateControl_update ? _GEN_1709 : _GEN_1741; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1774 = updateLogic_io_cacheUpdateControl_update ? _GEN_1710 : _GEN_1742; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1775 = updateLogic_io_cacheUpdateControl_update ? _GEN_1711 : _GEN_1743; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1776 = updateLogic_io_cacheUpdateControl_update ? _GEN_1712 : _GEN_1744; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1777 = updateLogic_io_cacheUpdateControl_update ? _GEN_1713 : _GEN_1745; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1778 = updateLogic_io_cacheUpdateControl_update ? _GEN_1714 : _GEN_1746; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1779 = updateLogic_io_cacheUpdateControl_update ? _GEN_1715 : _GEN_1747; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1780 = updateLogic_io_cacheUpdateControl_update ? _GEN_1716 : _GEN_1748; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1781 = updateLogic_io_cacheUpdateControl_update ? _GEN_1717 : _GEN_1749; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1782 = updateLogic_io_cacheUpdateControl_update ? _GEN_1718 : _GEN_1750; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1783 = updateLogic_io_cacheUpdateControl_update ? _GEN_1719 : _GEN_1751; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1784 = updateLogic_io_cacheUpdateControl_update ? _GEN_1720 : _GEN_1752; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1785 = updateLogic_io_cacheUpdateControl_update ? _GEN_1721 : _GEN_1753; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1786 = updateLogic_io_cacheUpdateControl_update ? _GEN_1722 : _GEN_1754; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1787 = updateLogic_io_cacheUpdateControl_update ? _GEN_1723 : _GEN_1755; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1788 = updateLogic_io_cacheUpdateControl_update ? _GEN_1724 : _GEN_1756; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1789 = updateLogic_io_cacheUpdateControl_update ? _GEN_1725 : _GEN_1757; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1790 = updateLogic_io_cacheUpdateControl_update ? _GEN_1726 : _GEN_1758; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1791 = updateLogic_io_cacheUpdateControl_update ? _GEN_1727 : _GEN_1759; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1792 = updateLogic_io_cacheUpdateControl_update ? _GEN_1728 : _GEN_1760; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1793 = updateLogic_io_cacheUpdateControl_update ? _GEN_1729 : _GEN_1761; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1794 = updateLogic_io_cacheUpdateControl_update ? _GEN_1730 : _GEN_1762; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1795 = updateLogic_io_cacheUpdateControl_update ? _GEN_1731 : _GEN_1763; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1796 = updateLogic_io_cacheUpdateControl_update ? _GEN_1732 : _GEN_1764; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1797 = updateLogic_io_cacheUpdateControl_update ? _GEN_1733 : _GEN_1765; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1798 = updateLogic_io_cacheUpdateControl_update ? _GEN_1734 : _GEN_1766; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1799 = updateLogic_io_cacheUpdateControl_update ? _GEN_1735 : _GEN_1767; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_1832 = _T_5 ? _GEN_1768 : REG_5_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1833 = _T_5 ? _GEN_1769 : REG_5_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1834 = _T_5 ? _GEN_1770 : REG_5_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1835 = _T_5 ? _GEN_1771 : REG_5_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1836 = _T_5 ? _GEN_1772 : REG_5_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1837 = _T_5 ? _GEN_1773 : REG_5_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1838 = _T_5 ? _GEN_1774 : REG_5_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1839 = _T_5 ? _GEN_1775 : REG_5_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1840 = _T_5 ? _GEN_1776 : REG_5_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1841 = _T_5 ? _GEN_1777 : REG_5_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1842 = _T_5 ? _GEN_1778 : REG_5_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1843 = _T_5 ? _GEN_1779 : REG_5_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1844 = _T_5 ? _GEN_1780 : REG_5_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1845 = _T_5 ? _GEN_1781 : REG_5_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1846 = _T_5 ? _GEN_1782 : REG_5_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1847 = _T_5 ? _GEN_1783 : REG_5_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1848 = _T_5 ? _GEN_1784 : REG_5_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1849 = _T_5 ? _GEN_1785 : REG_5_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1850 = _T_5 ? _GEN_1786 : REG_5_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1851 = _T_5 ? _GEN_1787 : REG_5_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1852 = _T_5 ? _GEN_1788 : REG_5_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1853 = _T_5 ? _GEN_1789 : REG_5_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1854 = _T_5 ? _GEN_1790 : REG_5_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1855 = _T_5 ? _GEN_1791 : REG_5_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1856 = _T_5 ? _GEN_1792 : REG_5_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1857 = _T_5 ? _GEN_1793 : REG_5_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1858 = _T_5 ? _GEN_1794 : REG_5_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1859 = _T_5 ? _GEN_1795 : REG_5_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1860 = _T_5 ? _GEN_1796 : REG_5_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1861 = _T_5 ? _GEN_1797 : REG_5_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1862 = _T_5 ? _GEN_1798 : REG_5_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1863 = _T_5 ? _GEN_1799 : REG_5_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_1864 = _GEN_2624 | _GEN_1832; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1865 = _GEN_2625 | _GEN_1833; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1866 = _GEN_2626 | _GEN_1834; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1867 = _GEN_2627 | _GEN_1835; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1868 = _GEN_2628 | _GEN_1836; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1869 = _GEN_2629 | _GEN_1837; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1870 = _GEN_2630 | _GEN_1838; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1871 = _GEN_2631 | _GEN_1839; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1872 = _GEN_2633 | _GEN_1840; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1873 = _GEN_2635 | _GEN_1841; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1874 = _GEN_2637 | _GEN_1842; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1875 = _GEN_2639 | _GEN_1843; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1876 = _GEN_2641 | _GEN_1844; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1877 = _GEN_2643 | _GEN_1845; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1878 = _GEN_2645 | _GEN_1846; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1879 = _GEN_2647 | _GEN_1847; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1880 = _GEN_2649 | _GEN_1848; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1881 = _GEN_2651 | _GEN_1849; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1882 = _GEN_2653 | _GEN_1850; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1883 = _GEN_2655 | _GEN_1851; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1884 = _GEN_2657 | _GEN_1852; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1885 = _GEN_2659 | _GEN_1853; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1886 = _GEN_2661 | _GEN_1854; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1887 = _GEN_2663 | _GEN_1855; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1888 = _GEN_2665 | _GEN_1856; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1889 = _GEN_2667 | _GEN_1857; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1890 = _GEN_2669 | _GEN_1858; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1891 = _GEN_2671 | _GEN_1859; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1892 = _GEN_2673 | _GEN_1860; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1893 = _GEN_2675 | _GEN_1861; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1894 = _GEN_2677 | _GEN_1862; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_1895 = _GEN_2679 | _GEN_1863; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_6 = MemBlock_6_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_1929 = 5'h1 == indexTagReg ? REG_14_1 : REG_14_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1930 = 5'h2 == indexTagReg ? REG_14_2 : _GEN_1929; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1931 = 5'h3 == indexTagReg ? REG_14_3 : _GEN_1930; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1932 = 5'h4 == indexTagReg ? REG_14_4 : _GEN_1931; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1933 = 5'h5 == indexTagReg ? REG_14_5 : _GEN_1932; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1934 = 5'h6 == indexTagReg ? REG_14_6 : _GEN_1933; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1935 = 5'h7 == indexTagReg ? REG_14_7 : _GEN_1934; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1936 = 5'h8 == indexTagReg ? REG_14_8 : _GEN_1935; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1937 = 5'h9 == indexTagReg ? REG_14_9 : _GEN_1936; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1938 = 5'ha == indexTagReg ? REG_14_10 : _GEN_1937; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1939 = 5'hb == indexTagReg ? REG_14_11 : _GEN_1938; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1940 = 5'hc == indexTagReg ? REG_14_12 : _GEN_1939; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1941 = 5'hd == indexTagReg ? REG_14_13 : _GEN_1940; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1942 = 5'he == indexTagReg ? REG_14_14 : _GEN_1941; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1943 = 5'hf == indexTagReg ? REG_14_15 : _GEN_1942; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1944 = 5'h10 == indexTagReg ? REG_14_16 : _GEN_1943; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1945 = 5'h11 == indexTagReg ? REG_14_17 : _GEN_1944; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1946 = 5'h12 == indexTagReg ? REG_14_18 : _GEN_1945; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1947 = 5'h13 == indexTagReg ? REG_14_19 : _GEN_1946; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1948 = 5'h14 == indexTagReg ? REG_14_20 : _GEN_1947; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1949 = 5'h15 == indexTagReg ? REG_14_21 : _GEN_1948; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1950 = 5'h16 == indexTagReg ? REG_14_22 : _GEN_1949; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1951 = 5'h17 == indexTagReg ? REG_14_23 : _GEN_1950; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1952 = 5'h18 == indexTagReg ? REG_14_24 : _GEN_1951; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1953 = 5'h19 == indexTagReg ? REG_14_25 : _GEN_1952; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1954 = 5'h1a == indexTagReg ? REG_14_26 : _GEN_1953; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1955 = 5'h1b == indexTagReg ? REG_14_27 : _GEN_1954; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1956 = 5'h1c == indexTagReg ? REG_14_28 : _GEN_1955; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1957 = 5'h1d == indexTagReg ? REG_14_29 : _GEN_1956; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1958 = 5'h1e == indexTagReg ? REG_14_30 : _GEN_1957; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_1959 = 5'h1f == indexTagReg ? REG_14_31 : _GEN_1958; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_6 = _GEN_1959 & tagTagReg == readTags_6; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_1961 = 5'h1 == indexTagReg ? REG_6_1 : REG_6_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1962 = 5'h2 == indexTagReg ? REG_6_2 : _GEN_1961; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1963 = 5'h3 == indexTagReg ? REG_6_3 : _GEN_1962; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1964 = 5'h4 == indexTagReg ? REG_6_4 : _GEN_1963; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1965 = 5'h5 == indexTagReg ? REG_6_5 : _GEN_1964; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1966 = 5'h6 == indexTagReg ? REG_6_6 : _GEN_1965; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1967 = 5'h7 == indexTagReg ? REG_6_7 : _GEN_1966; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1968 = 5'h8 == indexTagReg ? REG_6_8 : _GEN_1967; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1969 = 5'h9 == indexTagReg ? REG_6_9 : _GEN_1968; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1970 = 5'ha == indexTagReg ? REG_6_10 : _GEN_1969; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1971 = 5'hb == indexTagReg ? REG_6_11 : _GEN_1970; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1972 = 5'hc == indexTagReg ? REG_6_12 : _GEN_1971; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1973 = 5'hd == indexTagReg ? REG_6_13 : _GEN_1972; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1974 = 5'he == indexTagReg ? REG_6_14 : _GEN_1973; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1975 = 5'hf == indexTagReg ? REG_6_15 : _GEN_1974; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1976 = 5'h10 == indexTagReg ? REG_6_16 : _GEN_1975; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1977 = 5'h11 == indexTagReg ? REG_6_17 : _GEN_1976; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1978 = 5'h12 == indexTagReg ? REG_6_18 : _GEN_1977; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1979 = 5'h13 == indexTagReg ? REG_6_19 : _GEN_1978; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1980 = 5'h14 == indexTagReg ? REG_6_20 : _GEN_1979; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1981 = 5'h15 == indexTagReg ? REG_6_21 : _GEN_1980; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1982 = 5'h16 == indexTagReg ? REG_6_22 : _GEN_1981; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1983 = 5'h17 == indexTagReg ? REG_6_23 : _GEN_1982; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1984 = 5'h18 == indexTagReg ? REG_6_24 : _GEN_1983; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1985 = 5'h19 == indexTagReg ? REG_6_25 : _GEN_1984; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1986 = 5'h1a == indexTagReg ? REG_6_26 : _GEN_1985; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1987 = 5'h1b == indexTagReg ? REG_6_27 : _GEN_1986; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1988 = 5'h1c == indexTagReg ? REG_6_28 : _GEN_1987; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1989 = 5'h1d == indexTagReg ? REG_6_29 : _GEN_1988; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_1992 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_14_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1993 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_14_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1994 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_14_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1995 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_14_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1996 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_14_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1997 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_14_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1998 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_14_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_1999 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_14_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2000 = 4'h8 == _GEN_2632 | REG_14_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2001 = 4'h9 == _GEN_2632 | REG_14_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2002 = 4'ha == _GEN_2632 | REG_14_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2003 = 4'hb == _GEN_2632 | REG_14_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2004 = 4'hc == _GEN_2632 | REG_14_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2005 = 4'hd == _GEN_2632 | REG_14_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2006 = 4'he == _GEN_2632 | REG_14_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2007 = 4'hf == _GEN_2632 | REG_14_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2008 = 5'h10 == _GEN_2648 | REG_14_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2009 = 5'h11 == _GEN_2648 | REG_14_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2010 = 5'h12 == _GEN_2648 | REG_14_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2011 = 5'h13 == _GEN_2648 | REG_14_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2012 = 5'h14 == _GEN_2648 | REG_14_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2013 = 5'h15 == _GEN_2648 | REG_14_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2014 = 5'h16 == _GEN_2648 | REG_14_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2015 = 5'h17 == _GEN_2648 | REG_14_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2016 = 5'h18 == _GEN_2648 | REG_14_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2017 = 5'h19 == _GEN_2648 | REG_14_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2018 = 5'h1a == _GEN_2648 | REG_14_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2019 = 5'h1b == _GEN_2648 | REG_14_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2020 = 5'h1c == _GEN_2648 | REG_14_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2021 = 5'h1d == _GEN_2648 | REG_14_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2022 = 5'h1e == _GEN_2648 | REG_14_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2023 = 5'h1f == _GEN_2648 | REG_14_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2024 = _GEN_2624 | REG_6_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2025 = _GEN_2625 | REG_6_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2026 = _GEN_2626 | REG_6_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2027 = _GEN_2627 | REG_6_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2028 = _GEN_2628 | REG_6_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2029 = _GEN_2629 | REG_6_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2030 = _GEN_2630 | REG_6_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2031 = _GEN_2631 | REG_6_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2032 = _GEN_2633 | REG_6_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2033 = _GEN_2635 | REG_6_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2034 = _GEN_2637 | REG_6_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2035 = _GEN_2639 | REG_6_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2036 = _GEN_2641 | REG_6_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2037 = _GEN_2643 | REG_6_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2038 = _GEN_2645 | REG_6_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2039 = _GEN_2647 | REG_6_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2040 = _GEN_2649 | REG_6_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2041 = _GEN_2651 | REG_6_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2042 = _GEN_2653 | REG_6_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2043 = _GEN_2655 | REG_6_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2044 = _GEN_2657 | REG_6_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2045 = _GEN_2659 | REG_6_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2046 = _GEN_2661 | REG_6_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2047 = _GEN_2663 | REG_6_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2048 = _GEN_2665 | REG_6_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2049 = _GEN_2667 | REG_6_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2050 = _GEN_2669 | REG_6_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2051 = _GEN_2671 | REG_6_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2052 = _GEN_2673 | REG_6_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2053 = _GEN_2675 | REG_6_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2054 = _GEN_2677 | REG_6_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2055 = _GEN_2679 | REG_6_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2056 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2057 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2058 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2059 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2060 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2061 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2062 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2063 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_6_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2064 = 4'h8 == _GEN_2632 ? 1'h0 : REG_6_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2065 = 4'h9 == _GEN_2632 ? 1'h0 : REG_6_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2066 = 4'ha == _GEN_2632 ? 1'h0 : REG_6_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2067 = 4'hb == _GEN_2632 ? 1'h0 : REG_6_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2068 = 4'hc == _GEN_2632 ? 1'h0 : REG_6_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2069 = 4'hd == _GEN_2632 ? 1'h0 : REG_6_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2070 = 4'he == _GEN_2632 ? 1'h0 : REG_6_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2071 = 4'hf == _GEN_2632 ? 1'h0 : REG_6_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2072 = 5'h10 == _GEN_2648 ? 1'h0 : REG_6_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2073 = 5'h11 == _GEN_2648 ? 1'h0 : REG_6_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2074 = 5'h12 == _GEN_2648 ? 1'h0 : REG_6_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2075 = 5'h13 == _GEN_2648 ? 1'h0 : REG_6_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2076 = 5'h14 == _GEN_2648 ? 1'h0 : REG_6_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2077 = 5'h15 == _GEN_2648 ? 1'h0 : REG_6_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2078 = 5'h16 == _GEN_2648 ? 1'h0 : REG_6_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2079 = 5'h17 == _GEN_2648 ? 1'h0 : REG_6_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2080 = 5'h18 == _GEN_2648 ? 1'h0 : REG_6_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2081 = 5'h19 == _GEN_2648 ? 1'h0 : REG_6_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2082 = 5'h1a == _GEN_2648 ? 1'h0 : REG_6_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2083 = 5'h1b == _GEN_2648 ? 1'h0 : REG_6_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2084 = 5'h1c == _GEN_2648 ? 1'h0 : REG_6_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2085 = 5'h1d == _GEN_2648 ? 1'h0 : REG_6_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2086 = 5'h1e == _GEN_2648 ? 1'h0 : REG_6_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2087 = 5'h1f == _GEN_2648 ? 1'h0 : REG_6_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2088 = updateLogic_io_cacheUpdateControl_update ? _GEN_2024 : _GEN_2056; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2089 = updateLogic_io_cacheUpdateControl_update ? _GEN_2025 : _GEN_2057; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2090 = updateLogic_io_cacheUpdateControl_update ? _GEN_2026 : _GEN_2058; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2091 = updateLogic_io_cacheUpdateControl_update ? _GEN_2027 : _GEN_2059; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2092 = updateLogic_io_cacheUpdateControl_update ? _GEN_2028 : _GEN_2060; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2093 = updateLogic_io_cacheUpdateControl_update ? _GEN_2029 : _GEN_2061; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2094 = updateLogic_io_cacheUpdateControl_update ? _GEN_2030 : _GEN_2062; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2095 = updateLogic_io_cacheUpdateControl_update ? _GEN_2031 : _GEN_2063; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2096 = updateLogic_io_cacheUpdateControl_update ? _GEN_2032 : _GEN_2064; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2097 = updateLogic_io_cacheUpdateControl_update ? _GEN_2033 : _GEN_2065; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2098 = updateLogic_io_cacheUpdateControl_update ? _GEN_2034 : _GEN_2066; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2099 = updateLogic_io_cacheUpdateControl_update ? _GEN_2035 : _GEN_2067; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2100 = updateLogic_io_cacheUpdateControl_update ? _GEN_2036 : _GEN_2068; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2101 = updateLogic_io_cacheUpdateControl_update ? _GEN_2037 : _GEN_2069; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2102 = updateLogic_io_cacheUpdateControl_update ? _GEN_2038 : _GEN_2070; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2103 = updateLogic_io_cacheUpdateControl_update ? _GEN_2039 : _GEN_2071; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2104 = updateLogic_io_cacheUpdateControl_update ? _GEN_2040 : _GEN_2072; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2105 = updateLogic_io_cacheUpdateControl_update ? _GEN_2041 : _GEN_2073; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2106 = updateLogic_io_cacheUpdateControl_update ? _GEN_2042 : _GEN_2074; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2107 = updateLogic_io_cacheUpdateControl_update ? _GEN_2043 : _GEN_2075; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2108 = updateLogic_io_cacheUpdateControl_update ? _GEN_2044 : _GEN_2076; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2109 = updateLogic_io_cacheUpdateControl_update ? _GEN_2045 : _GEN_2077; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2110 = updateLogic_io_cacheUpdateControl_update ? _GEN_2046 : _GEN_2078; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2111 = updateLogic_io_cacheUpdateControl_update ? _GEN_2047 : _GEN_2079; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2112 = updateLogic_io_cacheUpdateControl_update ? _GEN_2048 : _GEN_2080; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2113 = updateLogic_io_cacheUpdateControl_update ? _GEN_2049 : _GEN_2081; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2114 = updateLogic_io_cacheUpdateControl_update ? _GEN_2050 : _GEN_2082; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2115 = updateLogic_io_cacheUpdateControl_update ? _GEN_2051 : _GEN_2083; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2116 = updateLogic_io_cacheUpdateControl_update ? _GEN_2052 : _GEN_2084; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2117 = updateLogic_io_cacheUpdateControl_update ? _GEN_2053 : _GEN_2085; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2118 = updateLogic_io_cacheUpdateControl_update ? _GEN_2054 : _GEN_2086; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2119 = updateLogic_io_cacheUpdateControl_update ? _GEN_2055 : _GEN_2087; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2152 = _T_6 ? _GEN_2088 : REG_6_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2153 = _T_6 ? _GEN_2089 : REG_6_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2154 = _T_6 ? _GEN_2090 : REG_6_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2155 = _T_6 ? _GEN_2091 : REG_6_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2156 = _T_6 ? _GEN_2092 : REG_6_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2157 = _T_6 ? _GEN_2093 : REG_6_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2158 = _T_6 ? _GEN_2094 : REG_6_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2159 = _T_6 ? _GEN_2095 : REG_6_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2160 = _T_6 ? _GEN_2096 : REG_6_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2161 = _T_6 ? _GEN_2097 : REG_6_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2162 = _T_6 ? _GEN_2098 : REG_6_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2163 = _T_6 ? _GEN_2099 : REG_6_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2164 = _T_6 ? _GEN_2100 : REG_6_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2165 = _T_6 ? _GEN_2101 : REG_6_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2166 = _T_6 ? _GEN_2102 : REG_6_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2167 = _T_6 ? _GEN_2103 : REG_6_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2168 = _T_6 ? _GEN_2104 : REG_6_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2169 = _T_6 ? _GEN_2105 : REG_6_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2170 = _T_6 ? _GEN_2106 : REG_6_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2171 = _T_6 ? _GEN_2107 : REG_6_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2172 = _T_6 ? _GEN_2108 : REG_6_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2173 = _T_6 ? _GEN_2109 : REG_6_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2174 = _T_6 ? _GEN_2110 : REG_6_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2175 = _T_6 ? _GEN_2111 : REG_6_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2176 = _T_6 ? _GEN_2112 : REG_6_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2177 = _T_6 ? _GEN_2113 : REG_6_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2178 = _T_6 ? _GEN_2114 : REG_6_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2179 = _T_6 ? _GEN_2115 : REG_6_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2180 = _T_6 ? _GEN_2116 : REG_6_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2181 = _T_6 ? _GEN_2117 : REG_6_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2182 = _T_6 ? _GEN_2118 : REG_6_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2183 = _T_6 ? _GEN_2119 : REG_6_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2184 = _GEN_2624 | _GEN_2152; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2185 = _GEN_2625 | _GEN_2153; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2186 = _GEN_2626 | _GEN_2154; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2187 = _GEN_2627 | _GEN_2155; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2188 = _GEN_2628 | _GEN_2156; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2189 = _GEN_2629 | _GEN_2157; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2190 = _GEN_2630 | _GEN_2158; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2191 = _GEN_2631 | _GEN_2159; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2192 = _GEN_2633 | _GEN_2160; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2193 = _GEN_2635 | _GEN_2161; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2194 = _GEN_2637 | _GEN_2162; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2195 = _GEN_2639 | _GEN_2163; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2196 = _GEN_2641 | _GEN_2164; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2197 = _GEN_2643 | _GEN_2165; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2198 = _GEN_2645 | _GEN_2166; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2199 = _GEN_2647 | _GEN_2167; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2200 = _GEN_2649 | _GEN_2168; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2201 = _GEN_2651 | _GEN_2169; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2202 = _GEN_2653 | _GEN_2170; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2203 = _GEN_2655 | _GEN_2171; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2204 = _GEN_2657 | _GEN_2172; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2205 = _GEN_2659 | _GEN_2173; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2206 = _GEN_2661 | _GEN_2174; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2207 = _GEN_2663 | _GEN_2175; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2208 = _GEN_2665 | _GEN_2176; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2209 = _GEN_2667 | _GEN_2177; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2210 = _GEN_2669 | _GEN_2178; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2211 = _GEN_2671 | _GEN_2179; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2212 = _GEN_2673 | _GEN_2180; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2213 = _GEN_2675 | _GEN_2181; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2214 = _GEN_2677 | _GEN_2182; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2215 = _GEN_2679 | _GEN_2183; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire [3:0] readTags_7 = MemBlock_7_io_readData; // @[SharedPipelinedCache.scala 73:22 84:22]
  wire  _GEN_2249 = 5'h1 == indexTagReg ? REG_15_1 : REG_15_0; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2250 = 5'h2 == indexTagReg ? REG_15_2 : _GEN_2249; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2251 = 5'h3 == indexTagReg ? REG_15_3 : _GEN_2250; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2252 = 5'h4 == indexTagReg ? REG_15_4 : _GEN_2251; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2253 = 5'h5 == indexTagReg ? REG_15_5 : _GEN_2252; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2254 = 5'h6 == indexTagReg ? REG_15_6 : _GEN_2253; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2255 = 5'h7 == indexTagReg ? REG_15_7 : _GEN_2254; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2256 = 5'h8 == indexTagReg ? REG_15_8 : _GEN_2255; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2257 = 5'h9 == indexTagReg ? REG_15_9 : _GEN_2256; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2258 = 5'ha == indexTagReg ? REG_15_10 : _GEN_2257; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2259 = 5'hb == indexTagReg ? REG_15_11 : _GEN_2258; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2260 = 5'hc == indexTagReg ? REG_15_12 : _GEN_2259; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2261 = 5'hd == indexTagReg ? REG_15_13 : _GEN_2260; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2262 = 5'he == indexTagReg ? REG_15_14 : _GEN_2261; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2263 = 5'hf == indexTagReg ? REG_15_15 : _GEN_2262; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2264 = 5'h10 == indexTagReg ? REG_15_16 : _GEN_2263; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2265 = 5'h11 == indexTagReg ? REG_15_17 : _GEN_2264; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2266 = 5'h12 == indexTagReg ? REG_15_18 : _GEN_2265; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2267 = 5'h13 == indexTagReg ? REG_15_19 : _GEN_2266; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2268 = 5'h14 == indexTagReg ? REG_15_20 : _GEN_2267; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2269 = 5'h15 == indexTagReg ? REG_15_21 : _GEN_2268; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2270 = 5'h16 == indexTagReg ? REG_15_22 : _GEN_2269; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2271 = 5'h17 == indexTagReg ? REG_15_23 : _GEN_2270; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2272 = 5'h18 == indexTagReg ? REG_15_24 : _GEN_2271; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2273 = 5'h19 == indexTagReg ? REG_15_25 : _GEN_2272; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2274 = 5'h1a == indexTagReg ? REG_15_26 : _GEN_2273; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2275 = 5'h1b == indexTagReg ? REG_15_27 : _GEN_2274; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2276 = 5'h1c == indexTagReg ? REG_15_28 : _GEN_2275; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2277 = 5'h1d == indexTagReg ? REG_15_29 : _GEN_2276; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2278 = 5'h1e == indexTagReg ? REG_15_30 : _GEN_2277; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  _GEN_2279 = 5'h1f == indexTagReg ? REG_15_31 : _GEN_2278; // @[SharedPipelinedCache.scala 106:{52,52}]
  wire  hits_7 = _GEN_2279 & tagTagReg == readTags_7; // @[SharedPipelinedCache.scala 106:52]
  wire  _GEN_2281 = 5'h1 == indexTagReg ? REG_7_1 : REG_7_0; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2282 = 5'h2 == indexTagReg ? REG_7_2 : _GEN_2281; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2283 = 5'h3 == indexTagReg ? REG_7_3 : _GEN_2282; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2284 = 5'h4 == indexTagReg ? REG_7_4 : _GEN_2283; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2285 = 5'h5 == indexTagReg ? REG_7_5 : _GEN_2284; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2286 = 5'h6 == indexTagReg ? REG_7_6 : _GEN_2285; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2287 = 5'h7 == indexTagReg ? REG_7_7 : _GEN_2286; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2288 = 5'h8 == indexTagReg ? REG_7_8 : _GEN_2287; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2289 = 5'h9 == indexTagReg ? REG_7_9 : _GEN_2288; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2290 = 5'ha == indexTagReg ? REG_7_10 : _GEN_2289; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2291 = 5'hb == indexTagReg ? REG_7_11 : _GEN_2290; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2292 = 5'hc == indexTagReg ? REG_7_12 : _GEN_2291; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2293 = 5'hd == indexTagReg ? REG_7_13 : _GEN_2292; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2294 = 5'he == indexTagReg ? REG_7_14 : _GEN_2293; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2295 = 5'hf == indexTagReg ? REG_7_15 : _GEN_2294; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2296 = 5'h10 == indexTagReg ? REG_7_16 : _GEN_2295; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2297 = 5'h11 == indexTagReg ? REG_7_17 : _GEN_2296; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2298 = 5'h12 == indexTagReg ? REG_7_18 : _GEN_2297; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2299 = 5'h13 == indexTagReg ? REG_7_19 : _GEN_2298; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2300 = 5'h14 == indexTagReg ? REG_7_20 : _GEN_2299; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2301 = 5'h15 == indexTagReg ? REG_7_21 : _GEN_2300; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2302 = 5'h16 == indexTagReg ? REG_7_22 : _GEN_2301; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2303 = 5'h17 == indexTagReg ? REG_7_23 : _GEN_2302; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2304 = 5'h18 == indexTagReg ? REG_7_24 : _GEN_2303; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2305 = 5'h19 == indexTagReg ? REG_7_25 : _GEN_2304; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2306 = 5'h1a == indexTagReg ? REG_7_26 : _GEN_2305; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2307 = 5'h1b == indexTagReg ? REG_7_27 : _GEN_2306; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2308 = 5'h1c == indexTagReg ? REG_7_28 : _GEN_2307; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2309 = 5'h1d == indexTagReg ? REG_7_29 : _GEN_2308; // @[SharedPipelinedCache.scala 107:{19,19}]
  wire  _GEN_2312 = 3'h0 == updateLogic_io_cacheUpdateControl_index | REG_15_0; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2313 = 3'h1 == updateLogic_io_cacheUpdateControl_index | REG_15_1; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2314 = 3'h2 == updateLogic_io_cacheUpdateControl_index | REG_15_2; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2315 = 3'h3 == updateLogic_io_cacheUpdateControl_index | REG_15_3; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2316 = 3'h4 == updateLogic_io_cacheUpdateControl_index | REG_15_4; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2317 = 3'h5 == updateLogic_io_cacheUpdateControl_index | REG_15_5; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2318 = 3'h6 == updateLogic_io_cacheUpdateControl_index | REG_15_6; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2319 = 3'h7 == updateLogic_io_cacheUpdateControl_index | REG_15_7; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2320 = 4'h8 == _GEN_2632 | REG_15_8; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2321 = 4'h9 == _GEN_2632 | REG_15_9; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2322 = 4'ha == _GEN_2632 | REG_15_10; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2323 = 4'hb == _GEN_2632 | REG_15_11; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2324 = 4'hc == _GEN_2632 | REG_15_12; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2325 = 4'hd == _GEN_2632 | REG_15_13; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2326 = 4'he == _GEN_2632 | REG_15_14; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2327 = 4'hf == _GEN_2632 | REG_15_15; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2328 = 5'h10 == _GEN_2648 | REG_15_16; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2329 = 5'h11 == _GEN_2648 | REG_15_17; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2330 = 5'h12 == _GEN_2648 | REG_15_18; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2331 = 5'h13 == _GEN_2648 | REG_15_19; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2332 = 5'h14 == _GEN_2648 | REG_15_20; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2333 = 5'h15 == _GEN_2648 | REG_15_21; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2334 = 5'h16 == _GEN_2648 | REG_15_22; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2335 = 5'h17 == _GEN_2648 | REG_15_23; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2336 = 5'h18 == _GEN_2648 | REG_15_24; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2337 = 5'h19 == _GEN_2648 | REG_15_25; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2338 = 5'h1a == _GEN_2648 | REG_15_26; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2339 = 5'h1b == _GEN_2648 | REG_15_27; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2340 = 5'h1c == _GEN_2648 | REG_15_28; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2341 = 5'h1d == _GEN_2648 | REG_15_29; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2342 = 5'h1e == _GEN_2648 | REG_15_30; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2343 = 5'h1f == _GEN_2648 | REG_15_31; // @[SharedPipelinedCache.scala 113:{66,66} 99:44]
  wire  _GEN_2344 = _GEN_2624 | REG_7_0; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2345 = _GEN_2625 | REG_7_1; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2346 = _GEN_2626 | REG_7_2; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2347 = _GEN_2627 | REG_7_3; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2348 = _GEN_2628 | REG_7_4; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2349 = _GEN_2629 | REG_7_5; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2350 = _GEN_2630 | REG_7_6; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2351 = _GEN_2631 | REG_7_7; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2352 = _GEN_2633 | REG_7_8; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2353 = _GEN_2635 | REG_7_9; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2354 = _GEN_2637 | REG_7_10; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2355 = _GEN_2639 | REG_7_11; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2356 = _GEN_2641 | REG_7_12; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2357 = _GEN_2643 | REG_7_13; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2358 = _GEN_2645 | REG_7_14; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2359 = _GEN_2647 | REG_7_15; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2360 = _GEN_2649 | REG_7_16; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2361 = _GEN_2651 | REG_7_17; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2362 = _GEN_2653 | REG_7_18; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2363 = _GEN_2655 | REG_7_19; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2364 = _GEN_2657 | REG_7_20; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2365 = _GEN_2659 | REG_7_21; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2366 = _GEN_2661 | REG_7_22; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2367 = _GEN_2663 | REG_7_23; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2368 = _GEN_2665 | REG_7_24; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2369 = _GEN_2667 | REG_7_25; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2370 = _GEN_2669 | REG_7_26; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2371 = _GEN_2671 | REG_7_27; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2372 = _GEN_2673 | REG_7_28; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2373 = _GEN_2675 | REG_7_29; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2374 = _GEN_2677 | REG_7_30; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2375 = _GEN_2679 | REG_7_31; // @[SharedPipelinedCache.scala 116:{68,68} 98:44]
  wire  _GEN_2376 = 3'h0 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_0; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2377 = 3'h1 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_1; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2378 = 3'h2 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_2; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2379 = 3'h3 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_3; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2380 = 3'h4 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_4; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2381 = 3'h5 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_5; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2382 = 3'h6 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_6; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2383 = 3'h7 == updateLogic_io_cacheUpdateControl_index ? 1'h0 : REG_7_7; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2384 = 4'h8 == _GEN_2632 ? 1'h0 : REG_7_8; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2385 = 4'h9 == _GEN_2632 ? 1'h0 : REG_7_9; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2386 = 4'ha == _GEN_2632 ? 1'h0 : REG_7_10; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2387 = 4'hb == _GEN_2632 ? 1'h0 : REG_7_11; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2388 = 4'hc == _GEN_2632 ? 1'h0 : REG_7_12; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2389 = 4'hd == _GEN_2632 ? 1'h0 : REG_7_13; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2390 = 4'he == _GEN_2632 ? 1'h0 : REG_7_14; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2391 = 4'hf == _GEN_2632 ? 1'h0 : REG_7_15; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2392 = 5'h10 == _GEN_2648 ? 1'h0 : REG_7_16; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2393 = 5'h11 == _GEN_2648 ? 1'h0 : REG_7_17; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2394 = 5'h12 == _GEN_2648 ? 1'h0 : REG_7_18; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2395 = 5'h13 == _GEN_2648 ? 1'h0 : REG_7_19; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2396 = 5'h14 == _GEN_2648 ? 1'h0 : REG_7_20; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2397 = 5'h15 == _GEN_2648 ? 1'h0 : REG_7_21; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2398 = 5'h16 == _GEN_2648 ? 1'h0 : REG_7_22; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2399 = 5'h17 == _GEN_2648 ? 1'h0 : REG_7_23; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2400 = 5'h18 == _GEN_2648 ? 1'h0 : REG_7_24; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2401 = 5'h19 == _GEN_2648 ? 1'h0 : REG_7_25; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2402 = 5'h1a == _GEN_2648 ? 1'h0 : REG_7_26; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2403 = 5'h1b == _GEN_2648 ? 1'h0 : REG_7_27; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2404 = 5'h1c == _GEN_2648 ? 1'h0 : REG_7_28; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2405 = 5'h1d == _GEN_2648 ? 1'h0 : REG_7_29; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2406 = 5'h1e == _GEN_2648 ? 1'h0 : REG_7_30; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2407 = 5'h1f == _GEN_2648 ? 1'h0 : REG_7_31; // @[SharedPipelinedCache.scala 118:{68,68} 98:44]
  wire  _GEN_2408 = updateLogic_io_cacheUpdateControl_update ? _GEN_2344 : _GEN_2376; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2409 = updateLogic_io_cacheUpdateControl_update ? _GEN_2345 : _GEN_2377; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2410 = updateLogic_io_cacheUpdateControl_update ? _GEN_2346 : _GEN_2378; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2411 = updateLogic_io_cacheUpdateControl_update ? _GEN_2347 : _GEN_2379; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2412 = updateLogic_io_cacheUpdateControl_update ? _GEN_2348 : _GEN_2380; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2413 = updateLogic_io_cacheUpdateControl_update ? _GEN_2349 : _GEN_2381; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2414 = updateLogic_io_cacheUpdateControl_update ? _GEN_2350 : _GEN_2382; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2415 = updateLogic_io_cacheUpdateControl_update ? _GEN_2351 : _GEN_2383; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2416 = updateLogic_io_cacheUpdateControl_update ? _GEN_2352 : _GEN_2384; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2417 = updateLogic_io_cacheUpdateControl_update ? _GEN_2353 : _GEN_2385; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2418 = updateLogic_io_cacheUpdateControl_update ? _GEN_2354 : _GEN_2386; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2419 = updateLogic_io_cacheUpdateControl_update ? _GEN_2355 : _GEN_2387; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2420 = updateLogic_io_cacheUpdateControl_update ? _GEN_2356 : _GEN_2388; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2421 = updateLogic_io_cacheUpdateControl_update ? _GEN_2357 : _GEN_2389; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2422 = updateLogic_io_cacheUpdateControl_update ? _GEN_2358 : _GEN_2390; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2423 = updateLogic_io_cacheUpdateControl_update ? _GEN_2359 : _GEN_2391; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2424 = updateLogic_io_cacheUpdateControl_update ? _GEN_2360 : _GEN_2392; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2425 = updateLogic_io_cacheUpdateControl_update ? _GEN_2361 : _GEN_2393; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2426 = updateLogic_io_cacheUpdateControl_update ? _GEN_2362 : _GEN_2394; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2427 = updateLogic_io_cacheUpdateControl_update ? _GEN_2363 : _GEN_2395; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2428 = updateLogic_io_cacheUpdateControl_update ? _GEN_2364 : _GEN_2396; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2429 = updateLogic_io_cacheUpdateControl_update ? _GEN_2365 : _GEN_2397; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2430 = updateLogic_io_cacheUpdateControl_update ? _GEN_2366 : _GEN_2398; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2431 = updateLogic_io_cacheUpdateControl_update ? _GEN_2367 : _GEN_2399; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2432 = updateLogic_io_cacheUpdateControl_update ? _GEN_2368 : _GEN_2400; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2433 = updateLogic_io_cacheUpdateControl_update ? _GEN_2369 : _GEN_2401; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2434 = updateLogic_io_cacheUpdateControl_update ? _GEN_2370 : _GEN_2402; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2435 = updateLogic_io_cacheUpdateControl_update ? _GEN_2371 : _GEN_2403; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2436 = updateLogic_io_cacheUpdateControl_update ? _GEN_2372 : _GEN_2404; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2437 = updateLogic_io_cacheUpdateControl_update ? _GEN_2373 : _GEN_2405; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2438 = updateLogic_io_cacheUpdateControl_update ? _GEN_2374 : _GEN_2406; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2439 = updateLogic_io_cacheUpdateControl_update ? _GEN_2375 : _GEN_2407; // @[SharedPipelinedCache.scala 115:54]
  wire  _GEN_2472 = _T_7 ? _GEN_2408 : REG_7_0; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2473 = _T_7 ? _GEN_2409 : REG_7_1; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2474 = _T_7 ? _GEN_2410 : REG_7_2; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2475 = _T_7 ? _GEN_2411 : REG_7_3; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2476 = _T_7 ? _GEN_2412 : REG_7_4; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2477 = _T_7 ? _GEN_2413 : REG_7_5; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2478 = _T_7 ? _GEN_2414 : REG_7_6; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2479 = _T_7 ? _GEN_2415 : REG_7_7; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2480 = _T_7 ? _GEN_2416 : REG_7_8; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2481 = _T_7 ? _GEN_2417 : REG_7_9; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2482 = _T_7 ? _GEN_2418 : REG_7_10; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2483 = _T_7 ? _GEN_2419 : REG_7_11; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2484 = _T_7 ? _GEN_2420 : REG_7_12; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2485 = _T_7 ? _GEN_2421 : REG_7_13; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2486 = _T_7 ? _GEN_2422 : REG_7_14; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2487 = _T_7 ? _GEN_2423 : REG_7_15; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2488 = _T_7 ? _GEN_2424 : REG_7_16; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2489 = _T_7 ? _GEN_2425 : REG_7_17; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2490 = _T_7 ? _GEN_2426 : REG_7_18; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2491 = _T_7 ? _GEN_2427 : REG_7_19; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2492 = _T_7 ? _GEN_2428 : REG_7_20; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2493 = _T_7 ? _GEN_2429 : REG_7_21; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2494 = _T_7 ? _GEN_2430 : REG_7_22; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2495 = _T_7 ? _GEN_2431 : REG_7_23; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2496 = _T_7 ? _GEN_2432 : REG_7_24; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2497 = _T_7 ? _GEN_2433 : REG_7_25; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2498 = _T_7 ? _GEN_2434 : REG_7_26; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2499 = _T_7 ? _GEN_2435 : REG_7_27; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2500 = _T_7 ? _GEN_2436 : REG_7_28; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2501 = _T_7 ? _GEN_2437 : REG_7_29; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2502 = _T_7 ? _GEN_2438 : REG_7_30; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2503 = _T_7 ? _GEN_2439 : REG_7_31; // @[SharedPipelinedCache.scala 112:67 98:44]
  wire  _GEN_2504 = _GEN_2624 | _GEN_2472; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2505 = _GEN_2625 | _GEN_2473; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2506 = _GEN_2626 | _GEN_2474; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2507 = _GEN_2627 | _GEN_2475; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2508 = _GEN_2628 | _GEN_2476; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2509 = _GEN_2629 | _GEN_2477; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2510 = _GEN_2630 | _GEN_2478; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2511 = _GEN_2631 | _GEN_2479; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2512 = _GEN_2633 | _GEN_2480; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2513 = _GEN_2635 | _GEN_2481; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2514 = _GEN_2637 | _GEN_2482; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2515 = _GEN_2639 | _GEN_2483; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2516 = _GEN_2641 | _GEN_2484; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2517 = _GEN_2643 | _GEN_2485; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2518 = _GEN_2645 | _GEN_2486; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2519 = _GEN_2647 | _GEN_2487; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2520 = _GEN_2649 | _GEN_2488; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2521 = _GEN_2651 | _GEN_2489; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2522 = _GEN_2653 | _GEN_2490; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2523 = _GEN_2655 | _GEN_2491; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2524 = _GEN_2657 | _GEN_2492; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2525 = _GEN_2659 | _GEN_2493; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2526 = _GEN_2661 | _GEN_2494; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2527 = _GEN_2663 | _GEN_2495; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2528 = _GEN_2665 | _GEN_2496; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2529 = _GEN_2667 | _GEN_2497; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2530 = _GEN_2669 | _GEN_2498; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2531 = _GEN_2671 | _GEN_2499; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2532 = _GEN_2673 | _GEN_2500; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2533 = _GEN_2675 | _GEN_2501; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2534 = _GEN_2677 | _GEN_2502; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  _GEN_2535 = _GEN_2679 | _GEN_2503; // @[SharedPipelinedCache.scala 124:{66,66}]
  wire  hit = hits_0 | hits_1 | hits_2 | hits_3 | hits_4 | hits_5 | hits_6 | hits_7; // @[SharedPipelinedCache.scala 128:37]
  wire [2:0] _hitWay_T = hits_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _hitWay_T_1 = hits_5 ? 3'h5 : _hitWay_T; // @[Mux.scala 47:70]
  wire [2:0] _hitWay_T_2 = hits_4 ? 3'h4 : _hitWay_T_1; // @[Mux.scala 47:70]
  wire [2:0] _hitWay_T_3 = hits_3 ? 3'h3 : _hitWay_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hitWay_T_4 = hits_2 ? 3'h2 : _hitWay_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hitWay_T_5 = hits_1 ? 3'h1 : _hitWay_T_4; // @[Mux.scala 47:70]
  wire [2:0] hitWay = hits_0 ? 3'h0 : _hitWay_T_5; // @[Mux.scala 47:70]
  reg [1:0] coreIdRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg  reqValidRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg [1:0] reqIdRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg  reqRwRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg [127:0] wDataRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg  hitRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg [2:0] hitWayRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_0; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_1; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_2; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_3; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_4; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_5; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_6; // @[SharedPipelinedCache.scala 42:30]
  reg  dirtyRepReg_7; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_0; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_1; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_2; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_3; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_4; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_5; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_6; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] readTagsRepReg_7; // @[SharedPipelinedCache.scala 42:30]
  reg [1:0] blockRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg [4:0] indexRepReg; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] tagRepReg; // @[SharedPipelinedCache.scala 42:30]
  wire  previousMissesCheck_0 = missQueue_io_currentIndexes_0 == indexRepReg & missQueue_io_currentWays_0 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_0; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_1 = missQueue_io_currentIndexes_1 == indexRepReg & missQueue_io_currentWays_1 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_1; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_2 = missQueue_io_currentIndexes_2 == indexRepReg & missQueue_io_currentWays_2 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_2; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_3 = missQueue_io_currentIndexes_3 == indexRepReg & missQueue_io_currentWays_3 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_3; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_4 = missQueue_io_currentIndexes_4 == indexRepReg & missQueue_io_currentWays_4 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_4; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_5 = missQueue_io_currentIndexes_5 == indexRepReg & missQueue_io_currentWays_5 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_5; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_6 = missQueue_io_currentIndexes_6 == indexRepReg & missQueue_io_currentWays_6 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_6; // @[SharedPipelinedCache.scala 166:82]
  wire  previousMissesCheck_7 = missQueue_io_currentIndexes_7 == indexRepReg & missQueue_io_currentWays_7 ==
    io_repPol_replaceWay & missQueue_io_validMSHRs_7; // @[SharedPipelinedCache.scala 166:82]
  wire  isPreviousMiss = previousMissesCheck_0 | previousMissesCheck_1 | previousMissesCheck_2 | previousMissesCheck_3
     | previousMissesCheck_4 | previousMissesCheck_5 | previousMissesCheck_6 | previousMissesCheck_7; // @[SharedPipelinedCache.scala 169:63]
  reg [1:0] coreIdReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg  reqValidReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg [1:0] reqIdReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg  reqRwReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg [127:0] wDataReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg  hitReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg [2:0] hitWayReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg  isRepDirtyReadReg; // @[SharedPipelinedCache.scala 42:30]
  wire  _GEN_2604 = 3'h1 == io_repPol_replaceWay ? dirtyRepReg_1 : dirtyRepReg_0; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire  _GEN_2605 = 3'h2 == io_repPol_replaceWay ? dirtyRepReg_2 : _GEN_2604; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire  _GEN_2606 = 3'h3 == io_repPol_replaceWay ? dirtyRepReg_3 : _GEN_2605; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire  _GEN_2607 = 3'h4 == io_repPol_replaceWay ? dirtyRepReg_4 : _GEN_2606; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire  _GEN_2608 = 3'h5 == io_repPol_replaceWay ? dirtyRepReg_5 : _GEN_2607; // @[SharedPipelinedCache.scala 44:{19,19}]
  reg [3:0] dirtyTagReadReg; // @[SharedPipelinedCache.scala 42:30]
  wire [3:0] _GEN_2613 = 3'h1 == io_repPol_replaceWay ? readTagsRepReg_1 : readTagsRepReg_0; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire [3:0] _GEN_2614 = 3'h2 == io_repPol_replaceWay ? readTagsRepReg_2 : _GEN_2613; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire [3:0] _GEN_2615 = 3'h3 == io_repPol_replaceWay ? readTagsRepReg_3 : _GEN_2614; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire [3:0] _GEN_2616 = 3'h4 == io_repPol_replaceWay ? readTagsRepReg_4 : _GEN_2615; // @[SharedPipelinedCache.scala 44:{19,19}]
  wire [3:0] _GEN_2617 = 3'h5 == io_repPol_replaceWay ? readTagsRepReg_5 : _GEN_2616; // @[SharedPipelinedCache.scala 44:{19,19}]
  reg [1:0] blockReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg [4:0] indexReadReg; // @[SharedPipelinedCache.scala 42:30]
  reg [3:0] tagReadReg; // @[SharedPipelinedCache.scala 42:30]
  wire [255:0] wbQueue_io_pushEntry_wbData_lo = {dataMem_io_rData_1,dataMem_io_rData_0}; // @[SharedPipelinedCache.scala 222:51]
  wire [255:0] wbQueue_io_pushEntry_wbData_hi = {dataMem_io_rData_3,dataMem_io_rData_2}; // @[SharedPipelinedCache.scala 222:51]
  MissFifo missQueue ( // @[SharedPipelinedCache.scala 49:25]
    .clock(missQueue_clock),
    .reset(missQueue_reset),
    .io_push(missQueue_io_push),
    .io_pushEntry_rw(missQueue_io_pushEntry_rw),
    .io_pushEntry_reqId(missQueue_io_pushEntry_reqId),
    .io_pushEntry_coreId(missQueue_io_pushEntry_coreId),
    .io_pushEntry_wData(missQueue_io_pushEntry_wData),
    .io_pushEntry_replaceWay(missQueue_io_pushEntry_replaceWay),
    .io_pushEntry_tag(missQueue_io_pushEntry_tag),
    .io_pushEntry_index(missQueue_io_pushEntry_index),
    .io_pushEntry_blockOffset(missQueue_io_pushEntry_blockOffset),
    .io_pop(missQueue_io_pop),
    .io_popEntry_rw(missQueue_io_popEntry_rw),
    .io_popEntry_reqId(missQueue_io_popEntry_reqId),
    .io_popEntry_coreId(missQueue_io_popEntry_coreId),
    .io_popEntry_wData(missQueue_io_popEntry_wData),
    .io_popEntry_replaceWay(missQueue_io_popEntry_replaceWay),
    .io_popEntry_tag(missQueue_io_popEntry_tag),
    .io_popEntry_index(missQueue_io_popEntry_index),
    .io_popEntry_blockOffset(missQueue_io_popEntry_blockOffset),
    .io_currentIndexes_0(missQueue_io_currentIndexes_0),
    .io_currentIndexes_1(missQueue_io_currentIndexes_1),
    .io_currentIndexes_2(missQueue_io_currentIndexes_2),
    .io_currentIndexes_3(missQueue_io_currentIndexes_3),
    .io_currentIndexes_4(missQueue_io_currentIndexes_4),
    .io_currentIndexes_5(missQueue_io_currentIndexes_5),
    .io_currentIndexes_6(missQueue_io_currentIndexes_6),
    .io_currentIndexes_7(missQueue_io_currentIndexes_7),
    .io_currentWays_0(missQueue_io_currentWays_0),
    .io_currentWays_1(missQueue_io_currentWays_1),
    .io_currentWays_2(missQueue_io_currentWays_2),
    .io_currentWays_3(missQueue_io_currentWays_3),
    .io_currentWays_4(missQueue_io_currentWays_4),
    .io_currentWays_5(missQueue_io_currentWays_5),
    .io_currentWays_6(missQueue_io_currentWays_6),
    .io_currentWays_7(missQueue_io_currentWays_7),
    .io_validMSHRs_0(missQueue_io_validMSHRs_0),
    .io_validMSHRs_1(missQueue_io_validMSHRs_1),
    .io_validMSHRs_2(missQueue_io_validMSHRs_2),
    .io_validMSHRs_3(missQueue_io_validMSHRs_3),
    .io_validMSHRs_4(missQueue_io_validMSHRs_4),
    .io_validMSHRs_5(missQueue_io_validMSHRs_5),
    .io_validMSHRs_6(missQueue_io_validMSHRs_6),
    .io_validMSHRs_7(missQueue_io_validMSHRs_7),
    .io_full(missQueue_io_full),
    .io_empty(missQueue_io_empty)
  );
  UpdateUnit updateLogic ( // @[SharedPipelinedCache.scala 50:27]
    .io_readStage_valid(updateLogic_io_readStage_valid),
    .io_readStage_reqId(updateLogic_io_readStage_reqId),
    .io_readStage_coreId(updateLogic_io_readStage_coreId),
    .io_readStage_rw(updateLogic_io_readStage_rw),
    .io_readStage_wData(updateLogic_io_readStage_wData),
    .io_readStage_wWay(updateLogic_io_readStage_wWay),
    .io_readStage_tag(updateLogic_io_readStage_tag),
    .io_readStage_index(updateLogic_io_readStage_index),
    .io_readStage_blockOffset(updateLogic_io_readStage_blockOffset),
    .io_readStage_memReadData_0(updateLogic_io_readStage_memReadData_0),
    .io_readStage_memReadData_1(updateLogic_io_readStage_memReadData_1),
    .io_readStage_memReadData_2(updateLogic_io_readStage_memReadData_2),
    .io_readStage_memReadData_3(updateLogic_io_readStage_memReadData_3),
    .io_memoryInterface_valid(updateLogic_io_memoryInterface_valid),
    .io_memoryInterface_reqId(updateLogic_io_memoryInterface_reqId),
    .io_memoryInterface_coreId(updateLogic_io_memoryInterface_coreId),
    .io_memoryInterface_rw(updateLogic_io_memoryInterface_rw),
    .io_memoryInterface_wData(updateLogic_io_memoryInterface_wData),
    .io_memoryInterface_wWay(updateLogic_io_memoryInterface_wWay),
    .io_memoryInterface_responseStatus(updateLogic_io_memoryInterface_responseStatus),
    .io_memoryInterface_tag(updateLogic_io_memoryInterface_tag),
    .io_memoryInterface_index(updateLogic_io_memoryInterface_index),
    .io_memoryInterface_blockOffset(updateLogic_io_memoryInterface_blockOffset),
    .io_memoryInterface_memReadData_0(updateLogic_io_memoryInterface_memReadData_0),
    .io_memoryInterface_memReadData_1(updateLogic_io_memoryInterface_memReadData_1),
    .io_memoryInterface_memReadData_2(updateLogic_io_memoryInterface_memReadData_2),
    .io_memoryInterface_memReadData_3(updateLogic_io_memoryInterface_memReadData_3),
    .io_cacheUpdateControl_tag(updateLogic_io_cacheUpdateControl_tag),
    .io_cacheUpdateControl_index(updateLogic_io_cacheUpdateControl_index),
    .io_cacheUpdateControl_coreId(updateLogic_io_cacheUpdateControl_coreId),
    .io_cacheUpdateControl_way(updateLogic_io_cacheUpdateControl_way),
    .io_cacheUpdateControl_refill(updateLogic_io_cacheUpdateControl_refill),
    .io_cacheUpdateControl_update(updateLogic_io_cacheUpdateControl_update),
    .io_cacheUpdateControl_stall(updateLogic_io_cacheUpdateControl_stall),
    .io_cacheUpdateControl_memWriteData_0(updateLogic_io_cacheUpdateControl_memWriteData_0),
    .io_cacheUpdateControl_memWriteData_1(updateLogic_io_cacheUpdateControl_memWriteData_1),
    .io_cacheUpdateControl_memWriteData_2(updateLogic_io_cacheUpdateControl_memWriteData_2),
    .io_cacheUpdateControl_memWriteData_3(updateLogic_io_cacheUpdateControl_memWriteData_3),
    .io_cacheUpdateControl_wrEn(updateLogic_io_cacheUpdateControl_wrEn),
    .io_coreResp_reqId_valid(updateLogic_io_coreResp_reqId_valid),
    .io_coreResp_reqId_bits(updateLogic_io_coreResp_reqId_bits),
    .io_coreResp_rData(updateLogic_io_coreResp_rData),
    .io_coreResp_responseStatus(updateLogic_io_coreResp_responseStatus)
  );
  RequestArbiter arbiter ( // @[SharedPipelinedCache.scala 55:23]
    .clock(arbiter_clock),
    .io_ports_0_reqId_ready(arbiter_io_ports_0_reqId_ready),
    .io_ports_0_reqId_valid(arbiter_io_ports_0_reqId_valid),
    .io_ports_0_reqId_bits(arbiter_io_ports_0_reqId_bits),
    .io_ports_0_addr(arbiter_io_ports_0_addr),
    .io_ports_0_rw(arbiter_io_ports_0_rw),
    .io_ports_0_wData(arbiter_io_ports_0_wData),
    .io_ports_1_reqId_ready(arbiter_io_ports_1_reqId_ready),
    .io_ports_1_reqId_valid(arbiter_io_ports_1_reqId_valid),
    .io_ports_1_reqId_bits(arbiter_io_ports_1_reqId_bits),
    .io_ports_1_addr(arbiter_io_ports_1_addr),
    .io_ports_1_rw(arbiter_io_ports_1_rw),
    .io_ports_1_wData(arbiter_io_ports_1_wData),
    .io_ports_2_reqId_ready(arbiter_io_ports_2_reqId_ready),
    .io_ports_2_reqId_valid(arbiter_io_ports_2_reqId_valid),
    .io_ports_2_reqId_bits(arbiter_io_ports_2_reqId_bits),
    .io_ports_2_addr(arbiter_io_ports_2_addr),
    .io_ports_2_rw(arbiter_io_ports_2_rw),
    .io_ports_2_wData(arbiter_io_ports_2_wData),
    .io_ports_3_reqId_ready(arbiter_io_ports_3_reqId_ready),
    .io_ports_3_reqId_valid(arbiter_io_ports_3_reqId_valid),
    .io_ports_3_reqId_bits(arbiter_io_ports_3_reqId_bits),
    .io_ports_3_addr(arbiter_io_ports_3_addr),
    .io_ports_3_rw(arbiter_io_ports_3_rw),
    .io_ports_3_wData(arbiter_io_ports_3_wData),
    .io_out_reqId_ready(arbiter_io_out_reqId_ready),
    .io_out_reqId_valid(arbiter_io_out_reqId_valid),
    .io_out_reqId_bits(arbiter_io_out_reqId_bits),
    .io_out_addr(arbiter_io_out_addr),
    .io_out_rw(arbiter_io_out_rw),
    .io_out_wData(arbiter_io_out_wData),
    .io_chosen(arbiter_io_chosen)
  );
  MemBlock MemBlock ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_clock),
    .io_readAddr(MemBlock_io_readAddr),
    .io_writeAddr(MemBlock_io_writeAddr),
    .io_writeData(MemBlock_io_writeData),
    .io_wrEn(MemBlock_io_wrEn),
    .io_readData(MemBlock_io_readData)
  );
  MemBlock MemBlock_1 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_1_clock),
    .io_readAddr(MemBlock_1_io_readAddr),
    .io_writeAddr(MemBlock_1_io_writeAddr),
    .io_writeData(MemBlock_1_io_writeData),
    .io_wrEn(MemBlock_1_io_wrEn),
    .io_readData(MemBlock_1_io_readData)
  );
  MemBlock MemBlock_2 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_2_clock),
    .io_readAddr(MemBlock_2_io_readAddr),
    .io_writeAddr(MemBlock_2_io_writeAddr),
    .io_writeData(MemBlock_2_io_writeData),
    .io_wrEn(MemBlock_2_io_wrEn),
    .io_readData(MemBlock_2_io_readData)
  );
  MemBlock MemBlock_3 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_3_clock),
    .io_readAddr(MemBlock_3_io_readAddr),
    .io_writeAddr(MemBlock_3_io_writeAddr),
    .io_writeData(MemBlock_3_io_writeData),
    .io_wrEn(MemBlock_3_io_wrEn),
    .io_readData(MemBlock_3_io_readData)
  );
  MemBlock MemBlock_4 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_4_clock),
    .io_readAddr(MemBlock_4_io_readAddr),
    .io_writeAddr(MemBlock_4_io_writeAddr),
    .io_writeData(MemBlock_4_io_writeData),
    .io_wrEn(MemBlock_4_io_wrEn),
    .io_readData(MemBlock_4_io_readData)
  );
  MemBlock MemBlock_5 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_5_clock),
    .io_readAddr(MemBlock_5_io_readAddr),
    .io_writeAddr(MemBlock_5_io_writeAddr),
    .io_writeData(MemBlock_5_io_writeData),
    .io_wrEn(MemBlock_5_io_wrEn),
    .io_readData(MemBlock_5_io_readData)
  );
  MemBlock MemBlock_6 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_6_clock),
    .io_readAddr(MemBlock_6_io_readAddr),
    .io_writeAddr(MemBlock_6_io_writeAddr),
    .io_writeData(MemBlock_6_io_writeData),
    .io_wrEn(MemBlock_6_io_wrEn),
    .io_readData(MemBlock_6_io_readData)
  );
  MemBlock MemBlock_7 ( // @[SharedPipelinedCache.scala 72:40]
    .clock(MemBlock_7_clock),
    .io_readAddr(MemBlock_7_io_readAddr),
    .io_writeAddr(MemBlock_7_io_writeAddr),
    .io_writeData(MemBlock_7_io_writeData),
    .io_wrEn(MemBlock_7_io_wrEn),
    .io_readData(MemBlock_7_io_readData)
  );
  CacheMemory dataMem ( // @[SharedPipelinedCache.scala 194:23]
    .clock(dataMem_clock),
    .io_rIndex(dataMem_io_rIndex),
    .io_rWayIdx(dataMem_io_rWayIdx),
    .io_wrIndex(dataMem_io_wrIndex),
    .io_wrWayIdx(dataMem_io_wrWayIdx),
    .io_wrEn(dataMem_io_wrEn),
    .io_wrData_0(dataMem_io_wrData_0),
    .io_wrData_1(dataMem_io_wrData_1),
    .io_wrData_2(dataMem_io_wrData_2),
    .io_wrData_3(dataMem_io_wrData_3),
    .io_rData_0(dataMem_io_rData_0),
    .io_rData_1(dataMem_io_rData_1),
    .io_rData_2(dataMem_io_rData_2),
    .io_rData_3(dataMem_io_rData_3)
  );
  WriteBackFifo wbQueue ( // @[SharedPipelinedCache.scala 219:23]
    .clock(wbQueue_clock),
    .reset(wbQueue_reset),
    .io_push(wbQueue_io_push),
    .io_pop(wbQueue_io_pop),
    .io_pushEntry_tag(wbQueue_io_pushEntry_tag),
    .io_pushEntry_index(wbQueue_io_pushEntry_index),
    .io_pushEntry_wbData(wbQueue_io_pushEntry_wbData),
    .io_popEntry_tag(wbQueue_io_popEntry_tag),
    .io_popEntry_index(wbQueue_io_popEntry_index),
    .io_popEntry_wbData(wbQueue_io_popEntry_wbData),
    .io_empty(wbQueue_io_empty)
  );
  MemoryInterface memInterface ( // @[SharedPipelinedCache.scala 228:28]
    .clock(memInterface_clock),
    .reset(memInterface_reset),
    .io_missFifo_popEntry_rw(memInterface_io_missFifo_popEntry_rw),
    .io_missFifo_popEntry_reqId(memInterface_io_missFifo_popEntry_reqId),
    .io_missFifo_popEntry_coreId(memInterface_io_missFifo_popEntry_coreId),
    .io_missFifo_popEntry_wData(memInterface_io_missFifo_popEntry_wData),
    .io_missFifo_popEntry_replaceWay(memInterface_io_missFifo_popEntry_replaceWay),
    .io_missFifo_popEntry_tag(memInterface_io_missFifo_popEntry_tag),
    .io_missFifo_popEntry_index(memInterface_io_missFifo_popEntry_index),
    .io_missFifo_popEntry_blockOffset(memInterface_io_missFifo_popEntry_blockOffset),
    .io_missFifo_empty(memInterface_io_missFifo_empty),
    .io_missFifo_pop(memInterface_io_missFifo_pop),
    .io_wbFifo_popEntry_tag(memInterface_io_wbFifo_popEntry_tag),
    .io_wbFifo_popEntry_index(memInterface_io_wbFifo_popEntry_index),
    .io_wbFifo_popEntry_wbData(memInterface_io_wbFifo_popEntry_wbData),
    .io_wbFifo_empty(memInterface_io_wbFifo_empty),
    .io_wbFifo_pop(memInterface_io_wbFifo_pop),
    .io_updateLogic_valid(memInterface_io_updateLogic_valid),
    .io_updateLogic_reqId(memInterface_io_updateLogic_reqId),
    .io_updateLogic_coreId(memInterface_io_updateLogic_coreId),
    .io_updateLogic_rw(memInterface_io_updateLogic_rw),
    .io_updateLogic_wData(memInterface_io_updateLogic_wData),
    .io_updateLogic_wWay(memInterface_io_updateLogic_wWay),
    .io_updateLogic_responseStatus(memInterface_io_updateLogic_responseStatus),
    .io_updateLogic_tag(memInterface_io_updateLogic_tag),
    .io_updateLogic_index(memInterface_io_updateLogic_index),
    .io_updateLogic_blockOffset(memInterface_io_updateLogic_blockOffset),
    .io_updateLogic_memReadData_0(memInterface_io_updateLogic_memReadData_0),
    .io_updateLogic_memReadData_1(memInterface_io_updateLogic_memReadData_1),
    .io_updateLogic_memReadData_2(memInterface_io_updateLogic_memReadData_2),
    .io_updateLogic_memReadData_3(memInterface_io_updateLogic_memReadData_3),
    .io_memController_rChannel_rAddr_ready(memInterface_io_memController_rChannel_rAddr_ready),
    .io_memController_rChannel_rAddr_valid(memInterface_io_memController_rChannel_rAddr_valid),
    .io_memController_rChannel_rAddr_bits(memInterface_io_memController_rChannel_rAddr_bits),
    .io_memController_rChannel_rData_ready(memInterface_io_memController_rChannel_rData_ready),
    .io_memController_rChannel_rData_valid(memInterface_io_memController_rChannel_rData_valid),
    .io_memController_rChannel_rData_bits(memInterface_io_memController_rChannel_rData_bits),
    .io_memController_rChannel_rLast(memInterface_io_memController_rChannel_rLast),
    .io_memController_wChannel_wAddr_ready(memInterface_io_memController_wChannel_wAddr_ready),
    .io_memController_wChannel_wAddr_valid(memInterface_io_memController_wChannel_wAddr_valid),
    .io_memController_wChannel_wAddr_bits(memInterface_io_memController_wChannel_wAddr_bits),
    .io_memController_wChannel_wData_ready(memInterface_io_memController_wChannel_wData_ready),
    .io_memController_wChannel_wData_valid(memInterface_io_memController_wChannel_wData_valid),
    .io_memController_wChannel_wData_bits(memInterface_io_memController_wChannel_wData_bits),
    .io_memController_wChannel_wLast(memInterface_io_memController_wChannel_wLast)
  );
  assign io_cache_coreReqs_0_reqId_ready = arbiter_io_ports_0_reqId_ready; // @[SharedPipelinedCache.scala 61:37]
  assign io_cache_coreReqs_1_reqId_ready = arbiter_io_ports_1_reqId_ready; // @[SharedPipelinedCache.scala 61:37]
  assign io_cache_coreReqs_2_reqId_ready = arbiter_io_ports_2_reqId_ready; // @[SharedPipelinedCache.scala 61:37]
  assign io_cache_coreReqs_3_reqId_ready = arbiter_io_ports_3_reqId_ready; // @[SharedPipelinedCache.scala 61:37]
  assign io_cache_coreResps_0_reqId_valid = updateLogic_io_cacheUpdateControl_coreId == 2'h0 &
    updateLogic_io_coreResp_reqId_valid; // @[SharedPipelinedCache.scala 257:105]
  assign io_cache_coreResps_0_reqId_bits = updateLogic_io_coreResp_reqId_bits; // @[SharedPipelinedCache.scala 258:44]
  assign io_cache_coreResps_0_rData = updateLogic_io_coreResp_rData; // @[SharedPipelinedCache.scala 259:39]
  assign io_cache_coreResps_0_responseStatus = updateLogic_io_coreResp_responseStatus; // @[SharedPipelinedCache.scala 260:48]
  assign io_cache_coreResps_1_reqId_valid = updateLogic_io_cacheUpdateControl_coreId == 2'h1 &
    updateLogic_io_coreResp_reqId_valid; // @[SharedPipelinedCache.scala 257:105]
  assign io_cache_coreResps_1_reqId_bits = updateLogic_io_coreResp_reqId_bits; // @[SharedPipelinedCache.scala 258:44]
  assign io_cache_coreResps_1_rData = updateLogic_io_coreResp_rData; // @[SharedPipelinedCache.scala 259:39]
  assign io_cache_coreResps_1_responseStatus = updateLogic_io_coreResp_responseStatus; // @[SharedPipelinedCache.scala 260:48]
  assign io_cache_coreResps_2_reqId_valid = updateLogic_io_cacheUpdateControl_coreId == 2'h2 &
    updateLogic_io_coreResp_reqId_valid; // @[SharedPipelinedCache.scala 257:105]
  assign io_cache_coreResps_2_reqId_bits = updateLogic_io_coreResp_reqId_bits; // @[SharedPipelinedCache.scala 258:44]
  assign io_cache_coreResps_2_rData = updateLogic_io_coreResp_rData; // @[SharedPipelinedCache.scala 259:39]
  assign io_cache_coreResps_2_responseStatus = updateLogic_io_coreResp_responseStatus; // @[SharedPipelinedCache.scala 260:48]
  assign io_cache_coreResps_3_reqId_valid = updateLogic_io_cacheUpdateControl_coreId == 2'h3 &
    updateLogic_io_coreResp_reqId_valid; // @[SharedPipelinedCache.scala 257:105]
  assign io_cache_coreResps_3_reqId_bits = updateLogic_io_coreResp_reqId_bits; // @[SharedPipelinedCache.scala 258:44]
  assign io_cache_coreResps_3_rData = updateLogic_io_coreResp_rData; // @[SharedPipelinedCache.scala 259:39]
  assign io_cache_coreResps_3_responseStatus = updateLogic_io_coreResp_responseStatus; // @[SharedPipelinedCache.scala 260:48]
  assign io_repPol_update_valid = reqValidTagReg; // @[SharedPipelinedCache.scala 131:26]
  assign io_repPol_update_bits = hit ? hitWay : io_repPol_replaceWay; // @[SharedPipelinedCache.scala 132:31]
  assign io_repPol_stall = updateLogic_io_cacheUpdateControl_stall; // @[SharedPipelinedCache.scala 134:19]
  assign io_repPol_setIdx = indexTagReg; // @[SharedPipelinedCache.scala 133:20]
  assign io_mem_rChannel_rAddr_valid = memInterface_io_memController_rChannel_rAddr_valid; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_rChannel_rAddr_bits = memInterface_io_memController_rChannel_rAddr_bits; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_rChannel_rData_ready = memInterface_io_memController_rChannel_rData_ready; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_wChannel_wAddr_valid = memInterface_io_memController_wChannel_wAddr_valid; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_wChannel_wAddr_bits = memInterface_io_memController_wChannel_wAddr_bits; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_wChannel_wData_valid = memInterface_io_memController_wChannel_wData_valid; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_wChannel_wData_bits = memInterface_io_memController_wChannel_wData_bits; // @[SharedPipelinedCache.scala 239:10]
  assign io_mem_wChannel_wLast = memInterface_io_memController_wChannel_wLast; // @[SharedPipelinedCache.scala 239:10]
  assign missQueue_clock = clock;
  assign missQueue_reset = reset;
  assign missQueue_io_push = isPreviousMiss | ~hitRepReg & reqValidRepReg; // @[SharedPipelinedCache.scala 177:23]
  assign missQueue_io_pushEntry_rw = reqRwRepReg; // @[SharedPipelinedCache.scala 185:29]
  assign missQueue_io_pushEntry_reqId = reqIdRepReg; // @[SharedPipelinedCache.scala 191:32]
  assign missQueue_io_pushEntry_coreId = coreIdRepReg; // @[SharedPipelinedCache.scala 192:33]
  assign missQueue_io_pushEntry_wData = wDataRepReg; // @[SharedPipelinedCache.scala 186:32]
  assign missQueue_io_pushEntry_replaceWay = io_repPol_replaceWay; // @[SharedPipelinedCache.scala 187:37]
  assign missQueue_io_pushEntry_tag = tagRepReg; // @[SharedPipelinedCache.scala 188:30]
  assign missQueue_io_pushEntry_index = indexRepReg; // @[SharedPipelinedCache.scala 189:32]
  assign missQueue_io_pushEntry_blockOffset = blockRepReg; // @[SharedPipelinedCache.scala 190:38]
  assign missQueue_io_pop = memInterface_io_missFifo_pop; // @[SharedPipelinedCache.scala 232:20]
  assign updateLogic_io_readStage_valid = reqValidReadReg & hitReadReg; // @[SharedPipelinedCache.scala 241:53]
  assign updateLogic_io_readStage_reqId = reqIdReadReg; // @[SharedPipelinedCache.scala 244:34]
  assign updateLogic_io_readStage_coreId = coreIdReadReg; // @[SharedPipelinedCache.scala 243:35]
  assign updateLogic_io_readStage_rw = reqRwReadReg; // @[SharedPipelinedCache.scala 242:31]
  assign updateLogic_io_readStage_wData = wDataReadReg; // @[SharedPipelinedCache.scala 245:34]
  assign updateLogic_io_readStage_wWay = hitWayReadReg; // @[SharedPipelinedCache.scala 246:33]
  assign updateLogic_io_readStage_tag = tagReadReg; // @[SharedPipelinedCache.scala 250:32]
  assign updateLogic_io_readStage_index = indexReadReg; // @[SharedPipelinedCache.scala 249:34]
  assign updateLogic_io_readStage_blockOffset = blockReadReg; // @[SharedPipelinedCache.scala 248:40]
  assign updateLogic_io_readStage_memReadData_0 = dataMem_io_rData_0; // @[SharedPipelinedCache.scala 251:40]
  assign updateLogic_io_readStage_memReadData_1 = dataMem_io_rData_1; // @[SharedPipelinedCache.scala 251:40]
  assign updateLogic_io_readStage_memReadData_2 = dataMem_io_rData_2; // @[SharedPipelinedCache.scala 251:40]
  assign updateLogic_io_readStage_memReadData_3 = dataMem_io_rData_3; // @[SharedPipelinedCache.scala 251:40]
  assign updateLogic_io_memoryInterface_valid = memInterface_io_updateLogic_valid; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_reqId = memInterface_io_updateLogic_reqId; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_coreId = memInterface_io_updateLogic_coreId; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_rw = memInterface_io_updateLogic_rw; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_wData = memInterface_io_updateLogic_wData; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_wWay = memInterface_io_updateLogic_wWay; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_responseStatus = memInterface_io_updateLogic_responseStatus; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_tag = memInterface_io_updateLogic_tag; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_index = memInterface_io_updateLogic_index; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_blockOffset = memInterface_io_updateLogic_blockOffset; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_memReadData_0 = memInterface_io_updateLogic_memReadData_0; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_memReadData_1 = memInterface_io_updateLogic_memReadData_1; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_memReadData_2 = memInterface_io_updateLogic_memReadData_2; // @[SharedPipelinedCache.scala 253:34]
  assign updateLogic_io_memoryInterface_memReadData_3 = memInterface_io_updateLogic_memReadData_3; // @[SharedPipelinedCache.scala 253:34]
  assign arbiter_clock = clock;
  assign arbiter_io_ports_0_reqId_valid = io_cache_coreReqs_0_reqId_valid; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_0_reqId_bits = io_cache_coreReqs_0_reqId_bits; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_0_addr = io_cache_coreReqs_0_addr; // @[SharedPipelinedCache.scala 62:36]
  assign arbiter_io_ports_0_rw = io_cache_coreReqs_0_rw; // @[SharedPipelinedCache.scala 63:34]
  assign arbiter_io_ports_0_wData = io_cache_coreReqs_0_wData; // @[SharedPipelinedCache.scala 64:37]
  assign arbiter_io_ports_1_reqId_valid = io_cache_coreReqs_1_reqId_valid; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_1_reqId_bits = io_cache_coreReqs_1_reqId_bits; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_1_addr = io_cache_coreReqs_1_addr; // @[SharedPipelinedCache.scala 62:36]
  assign arbiter_io_ports_1_rw = io_cache_coreReqs_1_rw; // @[SharedPipelinedCache.scala 63:34]
  assign arbiter_io_ports_1_wData = io_cache_coreReqs_1_wData; // @[SharedPipelinedCache.scala 64:37]
  assign arbiter_io_ports_2_reqId_valid = io_cache_coreReqs_2_reqId_valid; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_2_reqId_bits = io_cache_coreReqs_2_reqId_bits; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_2_addr = io_cache_coreReqs_2_addr; // @[SharedPipelinedCache.scala 62:36]
  assign arbiter_io_ports_2_rw = io_cache_coreReqs_2_rw; // @[SharedPipelinedCache.scala 63:34]
  assign arbiter_io_ports_2_wData = io_cache_coreReqs_2_wData; // @[SharedPipelinedCache.scala 64:37]
  assign arbiter_io_ports_3_reqId_valid = io_cache_coreReqs_3_reqId_valid; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_3_reqId_bits = io_cache_coreReqs_3_reqId_bits; // @[SharedPipelinedCache.scala 61:37]
  assign arbiter_io_ports_3_addr = io_cache_coreReqs_3_addr; // @[SharedPipelinedCache.scala 62:36]
  assign arbiter_io_ports_3_rw = io_cache_coreReqs_3_rw; // @[SharedPipelinedCache.scala 63:34]
  assign arbiter_io_ports_3_wData = io_cache_coreReqs_3_wData; // @[SharedPipelinedCache.scala 64:37]
  assign arbiter_io_out_reqId_ready = ~updateLogic_io_cacheUpdateControl_stall & ~missQueue_io_full; // @[SharedPipelinedCache.scala 56:30]
  assign MemBlock_clock = clock;
  assign MemBlock_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_1_clock = clock;
  assign MemBlock_1_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_1_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_1_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_1_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_1; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_2_clock = clock;
  assign MemBlock_2_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_2_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_2_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_2_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_2; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_3_clock = clock;
  assign MemBlock_3_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_3_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_3_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_3_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_3; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_4_clock = clock;
  assign MemBlock_4_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_4_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_4_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_4_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_4; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_5_clock = clock;
  assign MemBlock_5_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_5_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_5_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_5_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_5; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_6_clock = clock;
  assign MemBlock_6_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_6_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_6_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_6_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_6; // @[SharedPipelinedCache.scala 82:72]
  assign MemBlock_7_clock = clock;
  assign MemBlock_7_io_readAddr = arbiter_io_out_addr[10:6]; // @[SharedPipelinedCache.scala 69:34]
  assign MemBlock_7_io_writeAddr = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 81:33]
  assign MemBlock_7_io_writeData = updateLogic_io_cacheUpdateControl_tag; // @[SharedPipelinedCache.scala 80:33]
  assign MemBlock_7_io_wrEn = updateLogic_io_cacheUpdateControl_refill & isUpdateWay_7; // @[SharedPipelinedCache.scala 82:72]
  assign dataMem_clock = clock;
  assign dataMem_io_rIndex = indexRepReg; // @[SharedPipelinedCache.scala 196:21]
  assign dataMem_io_rWayIdx = hitRepReg ? hitWayRepReg : io_repPol_replaceWay; // @[SharedPipelinedCache.scala 197:28]
  assign dataMem_io_wrIndex = {{2'd0}, updateLogic_io_cacheUpdateControl_index}; // @[SharedPipelinedCache.scala 198:22]
  assign dataMem_io_wrWayIdx = updateLogic_io_cacheUpdateControl_way; // @[SharedPipelinedCache.scala 199:23]
  assign dataMem_io_wrEn = updateLogic_io_cacheUpdateControl_wrEn; // @[SharedPipelinedCache.scala 200:19]
  assign dataMem_io_wrData_0 = updateLogic_io_cacheUpdateControl_memWriteData_0; // @[SharedPipelinedCache.scala 201:21]
  assign dataMem_io_wrData_1 = updateLogic_io_cacheUpdateControl_memWriteData_1; // @[SharedPipelinedCache.scala 201:21]
  assign dataMem_io_wrData_2 = updateLogic_io_cacheUpdateControl_memWriteData_2; // @[SharedPipelinedCache.scala 201:21]
  assign dataMem_io_wrData_3 = updateLogic_io_cacheUpdateControl_memWriteData_3; // @[SharedPipelinedCache.scala 201:21]
  assign wbQueue_clock = clock;
  assign wbQueue_reset = reset;
  assign wbQueue_io_push = isRepDirtyReadReg & ~hitReadReg & reqValidReadReg; // @[SharedPipelinedCache.scala 221:55]
  assign wbQueue_io_pop = memInterface_io_wbFifo_pop; // @[SharedPipelinedCache.scala 236:18]
  assign wbQueue_io_pushEntry_tag = dirtyTagReadReg; // @[SharedPipelinedCache.scala 223:28]
  assign wbQueue_io_pushEntry_index = indexReadReg; // @[SharedPipelinedCache.scala 224:30]
  assign wbQueue_io_pushEntry_wbData = {wbQueue_io_pushEntry_wbData_hi,wbQueue_io_pushEntry_wbData_lo}; // @[SharedPipelinedCache.scala 222:51]
  assign memInterface_clock = clock;
  assign memInterface_reset = reset;
  assign memInterface_io_missFifo_popEntry_rw = missQueue_io_popEntry_rw; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_reqId = missQueue_io_popEntry_reqId; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_coreId = missQueue_io_popEntry_coreId; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_wData = missQueue_io_popEntry_wData; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_replaceWay = missQueue_io_popEntry_replaceWay; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_tag = missQueue_io_popEntry_tag; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_index = missQueue_io_popEntry_index; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_popEntry_blockOffset = missQueue_io_popEntry_blockOffset; // @[SharedPipelinedCache.scala 231:37]
  assign memInterface_io_missFifo_empty = missQueue_io_empty; // @[SharedPipelinedCache.scala 233:34]
  assign memInterface_io_wbFifo_popEntry_tag = wbQueue_io_popEntry_tag; // @[SharedPipelinedCache.scala 234:35]
  assign memInterface_io_wbFifo_popEntry_index = wbQueue_io_popEntry_index; // @[SharedPipelinedCache.scala 234:35]
  assign memInterface_io_wbFifo_popEntry_wbData = wbQueue_io_popEntry_wbData; // @[SharedPipelinedCache.scala 234:35]
  assign memInterface_io_wbFifo_empty = wbQueue_io_empty; // @[SharedPipelinedCache.scala 235:32]
  assign memInterface_io_memController_rChannel_rAddr_ready = io_mem_rChannel_rAddr_ready; // @[SharedPipelinedCache.scala 239:10]
  assign memInterface_io_memController_rChannel_rData_valid = io_mem_rChannel_rData_valid; // @[SharedPipelinedCache.scala 239:10]
  assign memInterface_io_memController_rChannel_rData_bits = io_mem_rChannel_rData_bits; // @[SharedPipelinedCache.scala 239:10]
  assign memInterface_io_memController_rChannel_rLast = io_mem_rChannel_rLast; // @[SharedPipelinedCache.scala 239:10]
  assign memInterface_io_memController_wChannel_wAddr_ready = io_mem_wChannel_wAddr_ready; // @[SharedPipelinedCache.scala 239:10]
  assign memInterface_io_memController_wChannel_wData_ready = io_mem_wChannel_wData_ready; // @[SharedPipelinedCache.scala 239:10]
  always @(posedge clock) begin
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      coreIdTagReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      coreIdTagReg <= arbiter_io_chosen; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqValidTagReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqValidTagReg <= _reqValidTagReg_T; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqIdTagReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqIdTagReg <= arbiter_io_out_reqId_bits; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqRwTagReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqRwTagReg <= arbiter_io_out_rw; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      wDataTagReg <= 128'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      wDataTagReg <= arbiter_io_out_wData; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      blockTagReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      blockTagReg <= blockOffset; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      indexTagReg <= 5'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      indexTagReg <= index; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      tagTagReg <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      tagTagReg <= tag; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__0 <= _GEN_264;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__0 <= _GEN_104;
      end else begin
        REG__0 <= _GEN_136;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__1 <= _GEN_265;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__1 <= _GEN_105;
      end else begin
        REG__1 <= _GEN_137;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__2 <= _GEN_266;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__2 <= _GEN_106;
      end else begin
        REG__2 <= _GEN_138;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__3 <= _GEN_267;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__3 <= _GEN_107;
      end else begin
        REG__3 <= _GEN_139;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__4 <= _GEN_268;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__4 <= _GEN_108;
      end else begin
        REG__4 <= _GEN_140;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__5 <= _GEN_269;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__5 <= _GEN_109;
      end else begin
        REG__5 <= _GEN_141;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__6 <= _GEN_270;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__6 <= _GEN_110;
      end else begin
        REG__6 <= _GEN_142;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__7 <= _GEN_271;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__7 <= _GEN_111;
      end else begin
        REG__7 <= _GEN_143;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__8 <= _GEN_272;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__8 <= _GEN_112;
      end else begin
        REG__8 <= _GEN_144;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__9 <= _GEN_273;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__9 <= _GEN_113;
      end else begin
        REG__9 <= _GEN_145;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__10 <= _GEN_274;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__10 <= _GEN_114;
      end else begin
        REG__10 <= _GEN_146;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__11 <= _GEN_275;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__11 <= _GEN_115;
      end else begin
        REG__11 <= _GEN_147;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__12 <= _GEN_276;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__12 <= _GEN_116;
      end else begin
        REG__12 <= _GEN_148;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__13 <= _GEN_277;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__13 <= _GEN_117;
      end else begin
        REG__13 <= _GEN_149;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__14 <= _GEN_278;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__14 <= _GEN_118;
      end else begin
        REG__14 <= _GEN_150;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__15 <= _GEN_279;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__15 <= _GEN_119;
      end else begin
        REG__15 <= _GEN_151;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__16 <= _GEN_280;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__16 <= _GEN_120;
      end else begin
        REG__16 <= _GEN_152;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__17 <= _GEN_281;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__17 <= _GEN_121;
      end else begin
        REG__17 <= _GEN_153;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__18 <= _GEN_282;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__18 <= _GEN_122;
      end else begin
        REG__18 <= _GEN_154;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__19 <= _GEN_283;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__19 <= _GEN_123;
      end else begin
        REG__19 <= _GEN_155;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__20 <= _GEN_284;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__20 <= _GEN_124;
      end else begin
        REG__20 <= _GEN_156;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__21 <= _GEN_285;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__21 <= _GEN_125;
      end else begin
        REG__21 <= _GEN_157;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__22 <= _GEN_286;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__22 <= _GEN_126;
      end else begin
        REG__22 <= _GEN_158;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__23 <= _GEN_287;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__23 <= _GEN_127;
      end else begin
        REG__23 <= _GEN_159;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__24 <= _GEN_288;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__24 <= _GEN_128;
      end else begin
        REG__24 <= _GEN_160;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__25 <= _GEN_289;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__25 <= _GEN_129;
      end else begin
        REG__25 <= _GEN_161;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__26 <= _GEN_290;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__26 <= _GEN_130;
      end else begin
        REG__26 <= _GEN_162;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__27 <= _GEN_291;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__27 <= _GEN_131;
      end else begin
        REG__27 <= _GEN_163;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__28 <= _GEN_292;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__28 <= _GEN_132;
      end else begin
        REG__28 <= _GEN_164;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__29 <= _GEN_293;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__29 <= _GEN_133;
      end else begin
        REG__29 <= _GEN_165;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__30 <= _GEN_294;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__30 <= _GEN_134;
      end else begin
        REG__30 <= _GEN_166;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG__31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG__31 <= _GEN_295;
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG__31 <= _GEN_135;
      end else begin
        REG__31 <= _GEN_167;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_0 <= _GEN_584;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_0 <= _GEN_424;
      end else begin
        REG_1_0 <= _GEN_456;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_1 <= _GEN_585;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_1 <= _GEN_425;
      end else begin
        REG_1_1 <= _GEN_457;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_2 <= _GEN_586;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_2 <= _GEN_426;
      end else begin
        REG_1_2 <= _GEN_458;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_3 <= _GEN_587;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_3 <= _GEN_427;
      end else begin
        REG_1_3 <= _GEN_459;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_4 <= _GEN_588;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_4 <= _GEN_428;
      end else begin
        REG_1_4 <= _GEN_460;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_5 <= _GEN_589;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_5 <= _GEN_429;
      end else begin
        REG_1_5 <= _GEN_461;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_6 <= _GEN_590;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_6 <= _GEN_430;
      end else begin
        REG_1_6 <= _GEN_462;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_7 <= _GEN_591;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_7 <= _GEN_431;
      end else begin
        REG_1_7 <= _GEN_463;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_8 <= _GEN_592;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_8 <= _GEN_432;
      end else begin
        REG_1_8 <= _GEN_464;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_9 <= _GEN_593;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_9 <= _GEN_433;
      end else begin
        REG_1_9 <= _GEN_465;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_10 <= _GEN_594;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_10 <= _GEN_434;
      end else begin
        REG_1_10 <= _GEN_466;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_11 <= _GEN_595;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_11 <= _GEN_435;
      end else begin
        REG_1_11 <= _GEN_467;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_12 <= _GEN_596;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_12 <= _GEN_436;
      end else begin
        REG_1_12 <= _GEN_468;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_13 <= _GEN_597;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_13 <= _GEN_437;
      end else begin
        REG_1_13 <= _GEN_469;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_14 <= _GEN_598;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_14 <= _GEN_438;
      end else begin
        REG_1_14 <= _GEN_470;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_15 <= _GEN_599;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_15 <= _GEN_439;
      end else begin
        REG_1_15 <= _GEN_471;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_16 <= _GEN_600;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_16 <= _GEN_440;
      end else begin
        REG_1_16 <= _GEN_472;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_17 <= _GEN_601;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_17 <= _GEN_441;
      end else begin
        REG_1_17 <= _GEN_473;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_18 <= _GEN_602;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_18 <= _GEN_442;
      end else begin
        REG_1_18 <= _GEN_474;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_19 <= _GEN_603;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_19 <= _GEN_443;
      end else begin
        REG_1_19 <= _GEN_475;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_20 <= _GEN_604;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_20 <= _GEN_444;
      end else begin
        REG_1_20 <= _GEN_476;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_21 <= _GEN_605;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_21 <= _GEN_445;
      end else begin
        REG_1_21 <= _GEN_477;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_22 <= _GEN_606;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_22 <= _GEN_446;
      end else begin
        REG_1_22 <= _GEN_478;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_23 <= _GEN_607;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_23 <= _GEN_447;
      end else begin
        REG_1_23 <= _GEN_479;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_24 <= _GEN_608;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_24 <= _GEN_448;
      end else begin
        REG_1_24 <= _GEN_480;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_25 <= _GEN_609;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_25 <= _GEN_449;
      end else begin
        REG_1_25 <= _GEN_481;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_26 <= _GEN_610;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_26 <= _GEN_450;
      end else begin
        REG_1_26 <= _GEN_482;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_27 <= _GEN_611;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_27 <= _GEN_451;
      end else begin
        REG_1_27 <= _GEN_483;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_28 <= _GEN_612;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_28 <= _GEN_452;
      end else begin
        REG_1_28 <= _GEN_484;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_29 <= _GEN_613;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_29 <= _GEN_453;
      end else begin
        REG_1_29 <= _GEN_485;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_30 <= _GEN_614;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_30 <= _GEN_454;
      end else begin
        REG_1_30 <= _GEN_486;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_1_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_1
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_1_31 <= _GEN_615;
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_1_31 <= _GEN_455;
      end else begin
        REG_1_31 <= _GEN_487;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_0 <= _GEN_904;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_0 <= _GEN_744;
      end else begin
        REG_2_0 <= _GEN_776;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_1 <= _GEN_905;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_1 <= _GEN_745;
      end else begin
        REG_2_1 <= _GEN_777;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_2 <= _GEN_906;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_2 <= _GEN_746;
      end else begin
        REG_2_2 <= _GEN_778;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_3 <= _GEN_907;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_3 <= _GEN_747;
      end else begin
        REG_2_3 <= _GEN_779;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_4 <= _GEN_908;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_4 <= _GEN_748;
      end else begin
        REG_2_4 <= _GEN_780;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_5 <= _GEN_909;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_5 <= _GEN_749;
      end else begin
        REG_2_5 <= _GEN_781;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_6 <= _GEN_910;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_6 <= _GEN_750;
      end else begin
        REG_2_6 <= _GEN_782;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_7 <= _GEN_911;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_7 <= _GEN_751;
      end else begin
        REG_2_7 <= _GEN_783;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_8 <= _GEN_912;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_8 <= _GEN_752;
      end else begin
        REG_2_8 <= _GEN_784;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_9 <= _GEN_913;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_9 <= _GEN_753;
      end else begin
        REG_2_9 <= _GEN_785;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_10 <= _GEN_914;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_10 <= _GEN_754;
      end else begin
        REG_2_10 <= _GEN_786;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_11 <= _GEN_915;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_11 <= _GEN_755;
      end else begin
        REG_2_11 <= _GEN_787;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_12 <= _GEN_916;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_12 <= _GEN_756;
      end else begin
        REG_2_12 <= _GEN_788;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_13 <= _GEN_917;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_13 <= _GEN_757;
      end else begin
        REG_2_13 <= _GEN_789;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_14 <= _GEN_918;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_14 <= _GEN_758;
      end else begin
        REG_2_14 <= _GEN_790;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_15 <= _GEN_919;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_15 <= _GEN_759;
      end else begin
        REG_2_15 <= _GEN_791;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_16 <= _GEN_920;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_16 <= _GEN_760;
      end else begin
        REG_2_16 <= _GEN_792;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_17 <= _GEN_921;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_17 <= _GEN_761;
      end else begin
        REG_2_17 <= _GEN_793;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_18 <= _GEN_922;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_18 <= _GEN_762;
      end else begin
        REG_2_18 <= _GEN_794;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_19 <= _GEN_923;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_19 <= _GEN_763;
      end else begin
        REG_2_19 <= _GEN_795;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_20 <= _GEN_924;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_20 <= _GEN_764;
      end else begin
        REG_2_20 <= _GEN_796;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_21 <= _GEN_925;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_21 <= _GEN_765;
      end else begin
        REG_2_21 <= _GEN_797;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_22 <= _GEN_926;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_22 <= _GEN_766;
      end else begin
        REG_2_22 <= _GEN_798;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_23 <= _GEN_927;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_23 <= _GEN_767;
      end else begin
        REG_2_23 <= _GEN_799;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_24 <= _GEN_928;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_24 <= _GEN_768;
      end else begin
        REG_2_24 <= _GEN_800;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_25 <= _GEN_929;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_25 <= _GEN_769;
      end else begin
        REG_2_25 <= _GEN_801;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_26 <= _GEN_930;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_26 <= _GEN_770;
      end else begin
        REG_2_26 <= _GEN_802;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_27 <= _GEN_931;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_27 <= _GEN_771;
      end else begin
        REG_2_27 <= _GEN_803;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_28 <= _GEN_932;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_28 <= _GEN_772;
      end else begin
        REG_2_28 <= _GEN_804;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_29 <= _GEN_933;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_29 <= _GEN_773;
      end else begin
        REG_2_29 <= _GEN_805;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_30 <= _GEN_934;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_30 <= _GEN_774;
      end else begin
        REG_2_30 <= _GEN_806;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_2_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_2
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_2_31 <= _GEN_935;
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_2_31 <= _GEN_775;
      end else begin
        REG_2_31 <= _GEN_807;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_0 <= _GEN_1224;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_0 <= _GEN_1064;
      end else begin
        REG_3_0 <= _GEN_1096;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_1 <= _GEN_1225;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_1 <= _GEN_1065;
      end else begin
        REG_3_1 <= _GEN_1097;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_2 <= _GEN_1226;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_2 <= _GEN_1066;
      end else begin
        REG_3_2 <= _GEN_1098;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_3 <= _GEN_1227;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_3 <= _GEN_1067;
      end else begin
        REG_3_3 <= _GEN_1099;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_4 <= _GEN_1228;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_4 <= _GEN_1068;
      end else begin
        REG_3_4 <= _GEN_1100;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_5 <= _GEN_1229;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_5 <= _GEN_1069;
      end else begin
        REG_3_5 <= _GEN_1101;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_6 <= _GEN_1230;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_6 <= _GEN_1070;
      end else begin
        REG_3_6 <= _GEN_1102;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_7 <= _GEN_1231;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_7 <= _GEN_1071;
      end else begin
        REG_3_7 <= _GEN_1103;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_8 <= _GEN_1232;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_8 <= _GEN_1072;
      end else begin
        REG_3_8 <= _GEN_1104;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_9 <= _GEN_1233;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_9 <= _GEN_1073;
      end else begin
        REG_3_9 <= _GEN_1105;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_10 <= _GEN_1234;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_10 <= _GEN_1074;
      end else begin
        REG_3_10 <= _GEN_1106;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_11 <= _GEN_1235;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_11 <= _GEN_1075;
      end else begin
        REG_3_11 <= _GEN_1107;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_12 <= _GEN_1236;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_12 <= _GEN_1076;
      end else begin
        REG_3_12 <= _GEN_1108;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_13 <= _GEN_1237;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_13 <= _GEN_1077;
      end else begin
        REG_3_13 <= _GEN_1109;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_14 <= _GEN_1238;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_14 <= _GEN_1078;
      end else begin
        REG_3_14 <= _GEN_1110;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_15 <= _GEN_1239;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_15 <= _GEN_1079;
      end else begin
        REG_3_15 <= _GEN_1111;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_16 <= _GEN_1240;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_16 <= _GEN_1080;
      end else begin
        REG_3_16 <= _GEN_1112;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_17 <= _GEN_1241;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_17 <= _GEN_1081;
      end else begin
        REG_3_17 <= _GEN_1113;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_18 <= _GEN_1242;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_18 <= _GEN_1082;
      end else begin
        REG_3_18 <= _GEN_1114;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_19 <= _GEN_1243;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_19 <= _GEN_1083;
      end else begin
        REG_3_19 <= _GEN_1115;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_20 <= _GEN_1244;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_20 <= _GEN_1084;
      end else begin
        REG_3_20 <= _GEN_1116;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_21 <= _GEN_1245;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_21 <= _GEN_1085;
      end else begin
        REG_3_21 <= _GEN_1117;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_22 <= _GEN_1246;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_22 <= _GEN_1086;
      end else begin
        REG_3_22 <= _GEN_1118;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_23 <= _GEN_1247;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_23 <= _GEN_1087;
      end else begin
        REG_3_23 <= _GEN_1119;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_24 <= _GEN_1248;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_24 <= _GEN_1088;
      end else begin
        REG_3_24 <= _GEN_1120;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_25 <= _GEN_1249;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_25 <= _GEN_1089;
      end else begin
        REG_3_25 <= _GEN_1121;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_26 <= _GEN_1250;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_26 <= _GEN_1090;
      end else begin
        REG_3_26 <= _GEN_1122;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_27 <= _GEN_1251;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_27 <= _GEN_1091;
      end else begin
        REG_3_27 <= _GEN_1123;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_28 <= _GEN_1252;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_28 <= _GEN_1092;
      end else begin
        REG_3_28 <= _GEN_1124;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_29 <= _GEN_1253;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_29 <= _GEN_1093;
      end else begin
        REG_3_29 <= _GEN_1125;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_30 <= _GEN_1254;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_30 <= _GEN_1094;
      end else begin
        REG_3_30 <= _GEN_1126;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_3_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_3
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_3_31 <= _GEN_1255;
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_3_31 <= _GEN_1095;
      end else begin
        REG_3_31 <= _GEN_1127;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_0 <= _GEN_1544;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_0 <= _GEN_1384;
      end else begin
        REG_4_0 <= _GEN_1416;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_1 <= _GEN_1545;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_1 <= _GEN_1385;
      end else begin
        REG_4_1 <= _GEN_1417;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_2 <= _GEN_1546;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_2 <= _GEN_1386;
      end else begin
        REG_4_2 <= _GEN_1418;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_3 <= _GEN_1547;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_3 <= _GEN_1387;
      end else begin
        REG_4_3 <= _GEN_1419;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_4 <= _GEN_1548;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_4 <= _GEN_1388;
      end else begin
        REG_4_4 <= _GEN_1420;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_5 <= _GEN_1549;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_5 <= _GEN_1389;
      end else begin
        REG_4_5 <= _GEN_1421;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_6 <= _GEN_1550;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_6 <= _GEN_1390;
      end else begin
        REG_4_6 <= _GEN_1422;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_7 <= _GEN_1551;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_7 <= _GEN_1391;
      end else begin
        REG_4_7 <= _GEN_1423;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_8 <= _GEN_1552;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_8 <= _GEN_1392;
      end else begin
        REG_4_8 <= _GEN_1424;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_9 <= _GEN_1553;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_9 <= _GEN_1393;
      end else begin
        REG_4_9 <= _GEN_1425;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_10 <= _GEN_1554;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_10 <= _GEN_1394;
      end else begin
        REG_4_10 <= _GEN_1426;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_11 <= _GEN_1555;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_11 <= _GEN_1395;
      end else begin
        REG_4_11 <= _GEN_1427;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_12 <= _GEN_1556;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_12 <= _GEN_1396;
      end else begin
        REG_4_12 <= _GEN_1428;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_13 <= _GEN_1557;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_13 <= _GEN_1397;
      end else begin
        REG_4_13 <= _GEN_1429;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_14 <= _GEN_1558;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_14 <= _GEN_1398;
      end else begin
        REG_4_14 <= _GEN_1430;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_15 <= _GEN_1559;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_15 <= _GEN_1399;
      end else begin
        REG_4_15 <= _GEN_1431;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_16 <= _GEN_1560;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_16 <= _GEN_1400;
      end else begin
        REG_4_16 <= _GEN_1432;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_17 <= _GEN_1561;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_17 <= _GEN_1401;
      end else begin
        REG_4_17 <= _GEN_1433;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_18 <= _GEN_1562;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_18 <= _GEN_1402;
      end else begin
        REG_4_18 <= _GEN_1434;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_19 <= _GEN_1563;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_19 <= _GEN_1403;
      end else begin
        REG_4_19 <= _GEN_1435;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_20 <= _GEN_1564;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_20 <= _GEN_1404;
      end else begin
        REG_4_20 <= _GEN_1436;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_21 <= _GEN_1565;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_21 <= _GEN_1405;
      end else begin
        REG_4_21 <= _GEN_1437;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_22 <= _GEN_1566;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_22 <= _GEN_1406;
      end else begin
        REG_4_22 <= _GEN_1438;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_23 <= _GEN_1567;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_23 <= _GEN_1407;
      end else begin
        REG_4_23 <= _GEN_1439;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_24 <= _GEN_1568;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_24 <= _GEN_1408;
      end else begin
        REG_4_24 <= _GEN_1440;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_25 <= _GEN_1569;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_25 <= _GEN_1409;
      end else begin
        REG_4_25 <= _GEN_1441;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_26 <= _GEN_1570;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_26 <= _GEN_1410;
      end else begin
        REG_4_26 <= _GEN_1442;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_27 <= _GEN_1571;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_27 <= _GEN_1411;
      end else begin
        REG_4_27 <= _GEN_1443;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_28 <= _GEN_1572;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_28 <= _GEN_1412;
      end else begin
        REG_4_28 <= _GEN_1444;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_29 <= _GEN_1573;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_29 <= _GEN_1413;
      end else begin
        REG_4_29 <= _GEN_1445;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_30 <= _GEN_1574;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_30 <= _GEN_1414;
      end else begin
        REG_4_30 <= _GEN_1446;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_4_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_4
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_4_31 <= _GEN_1575;
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_4_31 <= _GEN_1415;
      end else begin
        REG_4_31 <= _GEN_1447;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_0 <= _GEN_1864;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_0 <= _GEN_1704;
      end else begin
        REG_5_0 <= _GEN_1736;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_1 <= _GEN_1865;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_1 <= _GEN_1705;
      end else begin
        REG_5_1 <= _GEN_1737;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_2 <= _GEN_1866;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_2 <= _GEN_1706;
      end else begin
        REG_5_2 <= _GEN_1738;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_3 <= _GEN_1867;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_3 <= _GEN_1707;
      end else begin
        REG_5_3 <= _GEN_1739;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_4 <= _GEN_1868;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_4 <= _GEN_1708;
      end else begin
        REG_5_4 <= _GEN_1740;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_5 <= _GEN_1869;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_5 <= _GEN_1709;
      end else begin
        REG_5_5 <= _GEN_1741;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_6 <= _GEN_1870;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_6 <= _GEN_1710;
      end else begin
        REG_5_6 <= _GEN_1742;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_7 <= _GEN_1871;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_7 <= _GEN_1711;
      end else begin
        REG_5_7 <= _GEN_1743;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_8 <= _GEN_1872;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_8 <= _GEN_1712;
      end else begin
        REG_5_8 <= _GEN_1744;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_9 <= _GEN_1873;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_9 <= _GEN_1713;
      end else begin
        REG_5_9 <= _GEN_1745;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_10 <= _GEN_1874;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_10 <= _GEN_1714;
      end else begin
        REG_5_10 <= _GEN_1746;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_11 <= _GEN_1875;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_11 <= _GEN_1715;
      end else begin
        REG_5_11 <= _GEN_1747;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_12 <= _GEN_1876;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_12 <= _GEN_1716;
      end else begin
        REG_5_12 <= _GEN_1748;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_13 <= _GEN_1877;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_13 <= _GEN_1717;
      end else begin
        REG_5_13 <= _GEN_1749;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_14 <= _GEN_1878;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_14 <= _GEN_1718;
      end else begin
        REG_5_14 <= _GEN_1750;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_15 <= _GEN_1879;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_15 <= _GEN_1719;
      end else begin
        REG_5_15 <= _GEN_1751;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_16 <= _GEN_1880;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_16 <= _GEN_1720;
      end else begin
        REG_5_16 <= _GEN_1752;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_17 <= _GEN_1881;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_17 <= _GEN_1721;
      end else begin
        REG_5_17 <= _GEN_1753;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_18 <= _GEN_1882;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_18 <= _GEN_1722;
      end else begin
        REG_5_18 <= _GEN_1754;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_19 <= _GEN_1883;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_19 <= _GEN_1723;
      end else begin
        REG_5_19 <= _GEN_1755;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_20 <= _GEN_1884;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_20 <= _GEN_1724;
      end else begin
        REG_5_20 <= _GEN_1756;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_21 <= _GEN_1885;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_21 <= _GEN_1725;
      end else begin
        REG_5_21 <= _GEN_1757;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_22 <= _GEN_1886;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_22 <= _GEN_1726;
      end else begin
        REG_5_22 <= _GEN_1758;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_23 <= _GEN_1887;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_23 <= _GEN_1727;
      end else begin
        REG_5_23 <= _GEN_1759;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_24 <= _GEN_1888;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_24 <= _GEN_1728;
      end else begin
        REG_5_24 <= _GEN_1760;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_25 <= _GEN_1889;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_25 <= _GEN_1729;
      end else begin
        REG_5_25 <= _GEN_1761;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_26 <= _GEN_1890;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_26 <= _GEN_1730;
      end else begin
        REG_5_26 <= _GEN_1762;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_27 <= _GEN_1891;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_27 <= _GEN_1731;
      end else begin
        REG_5_27 <= _GEN_1763;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_28 <= _GEN_1892;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_28 <= _GEN_1732;
      end else begin
        REG_5_28 <= _GEN_1764;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_29 <= _GEN_1893;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_29 <= _GEN_1733;
      end else begin
        REG_5_29 <= _GEN_1765;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_30 <= _GEN_1894;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_30 <= _GEN_1734;
      end else begin
        REG_5_30 <= _GEN_1766;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_5_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_5
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_5_31 <= _GEN_1895;
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_5_31 <= _GEN_1735;
      end else begin
        REG_5_31 <= _GEN_1767;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_0 <= _GEN_2184;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_0 <= _GEN_2024;
      end else begin
        REG_6_0 <= _GEN_2056;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_1 <= _GEN_2185;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_1 <= _GEN_2025;
      end else begin
        REG_6_1 <= _GEN_2057;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_2 <= _GEN_2186;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_2 <= _GEN_2026;
      end else begin
        REG_6_2 <= _GEN_2058;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_3 <= _GEN_2187;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_3 <= _GEN_2027;
      end else begin
        REG_6_3 <= _GEN_2059;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_4 <= _GEN_2188;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_4 <= _GEN_2028;
      end else begin
        REG_6_4 <= _GEN_2060;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_5 <= _GEN_2189;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_5 <= _GEN_2029;
      end else begin
        REG_6_5 <= _GEN_2061;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_6 <= _GEN_2190;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_6 <= _GEN_2030;
      end else begin
        REG_6_6 <= _GEN_2062;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_7 <= _GEN_2191;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_7 <= _GEN_2031;
      end else begin
        REG_6_7 <= _GEN_2063;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_8 <= _GEN_2192;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_8 <= _GEN_2032;
      end else begin
        REG_6_8 <= _GEN_2064;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_9 <= _GEN_2193;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_9 <= _GEN_2033;
      end else begin
        REG_6_9 <= _GEN_2065;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_10 <= _GEN_2194;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_10 <= _GEN_2034;
      end else begin
        REG_6_10 <= _GEN_2066;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_11 <= _GEN_2195;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_11 <= _GEN_2035;
      end else begin
        REG_6_11 <= _GEN_2067;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_12 <= _GEN_2196;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_12 <= _GEN_2036;
      end else begin
        REG_6_12 <= _GEN_2068;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_13 <= _GEN_2197;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_13 <= _GEN_2037;
      end else begin
        REG_6_13 <= _GEN_2069;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_14 <= _GEN_2198;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_14 <= _GEN_2038;
      end else begin
        REG_6_14 <= _GEN_2070;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_15 <= _GEN_2199;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_15 <= _GEN_2039;
      end else begin
        REG_6_15 <= _GEN_2071;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_16 <= _GEN_2200;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_16 <= _GEN_2040;
      end else begin
        REG_6_16 <= _GEN_2072;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_17 <= _GEN_2201;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_17 <= _GEN_2041;
      end else begin
        REG_6_17 <= _GEN_2073;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_18 <= _GEN_2202;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_18 <= _GEN_2042;
      end else begin
        REG_6_18 <= _GEN_2074;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_19 <= _GEN_2203;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_19 <= _GEN_2043;
      end else begin
        REG_6_19 <= _GEN_2075;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_20 <= _GEN_2204;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_20 <= _GEN_2044;
      end else begin
        REG_6_20 <= _GEN_2076;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_21 <= _GEN_2205;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_21 <= _GEN_2045;
      end else begin
        REG_6_21 <= _GEN_2077;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_22 <= _GEN_2206;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_22 <= _GEN_2046;
      end else begin
        REG_6_22 <= _GEN_2078;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_23 <= _GEN_2207;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_23 <= _GEN_2047;
      end else begin
        REG_6_23 <= _GEN_2079;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_24 <= _GEN_2208;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_24 <= _GEN_2048;
      end else begin
        REG_6_24 <= _GEN_2080;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_25 <= _GEN_2209;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_25 <= _GEN_2049;
      end else begin
        REG_6_25 <= _GEN_2081;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_26 <= _GEN_2210;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_26 <= _GEN_2050;
      end else begin
        REG_6_26 <= _GEN_2082;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_27 <= _GEN_2211;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_27 <= _GEN_2051;
      end else begin
        REG_6_27 <= _GEN_2083;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_28 <= _GEN_2212;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_28 <= _GEN_2052;
      end else begin
        REG_6_28 <= _GEN_2084;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_29 <= _GEN_2213;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_29 <= _GEN_2053;
      end else begin
        REG_6_29 <= _GEN_2085;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_30 <= _GEN_2214;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_30 <= _GEN_2054;
      end else begin
        REG_6_30 <= _GEN_2086;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_6_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_6
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_6_31 <= _GEN_2215;
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_6_31 <= _GEN_2055;
      end else begin
        REG_6_31 <= _GEN_2087;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_0 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_0 <= _GEN_2504;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_0 <= _GEN_2344;
      end else begin
        REG_7_0 <= _GEN_2376;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_1 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_1 <= _GEN_2505;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_1 <= _GEN_2345;
      end else begin
        REG_7_1 <= _GEN_2377;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_2 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_2 <= _GEN_2506;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_2 <= _GEN_2346;
      end else begin
        REG_7_2 <= _GEN_2378;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_3 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_3 <= _GEN_2507;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_3 <= _GEN_2347;
      end else begin
        REG_7_3 <= _GEN_2379;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_4 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_4 <= _GEN_2508;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_4 <= _GEN_2348;
      end else begin
        REG_7_4 <= _GEN_2380;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_5 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_5 <= _GEN_2509;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_5 <= _GEN_2349;
      end else begin
        REG_7_5 <= _GEN_2381;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_6 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_6 <= _GEN_2510;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_6 <= _GEN_2350;
      end else begin
        REG_7_6 <= _GEN_2382;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_7 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_7 <= _GEN_2511;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_7 <= _GEN_2351;
      end else begin
        REG_7_7 <= _GEN_2383;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_8 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_8 <= _GEN_2512;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_8 <= _GEN_2352;
      end else begin
        REG_7_8 <= _GEN_2384;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_9 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_9 <= _GEN_2513;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_9 <= _GEN_2353;
      end else begin
        REG_7_9 <= _GEN_2385;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_10 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_10 <= _GEN_2514;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_10 <= _GEN_2354;
      end else begin
        REG_7_10 <= _GEN_2386;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_11 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_11 <= _GEN_2515;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_11 <= _GEN_2355;
      end else begin
        REG_7_11 <= _GEN_2387;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_12 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_12 <= _GEN_2516;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_12 <= _GEN_2356;
      end else begin
        REG_7_12 <= _GEN_2388;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_13 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_13 <= _GEN_2517;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_13 <= _GEN_2357;
      end else begin
        REG_7_13 <= _GEN_2389;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_14 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_14 <= _GEN_2518;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_14 <= _GEN_2358;
      end else begin
        REG_7_14 <= _GEN_2390;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_15 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_15 <= _GEN_2519;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_15 <= _GEN_2359;
      end else begin
        REG_7_15 <= _GEN_2391;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_16 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_16 <= _GEN_2520;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_16 <= _GEN_2360;
      end else begin
        REG_7_16 <= _GEN_2392;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_17 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_17 <= _GEN_2521;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_17 <= _GEN_2361;
      end else begin
        REG_7_17 <= _GEN_2393;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_18 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_18 <= _GEN_2522;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_18 <= _GEN_2362;
      end else begin
        REG_7_18 <= _GEN_2394;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_19 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_19 <= _GEN_2523;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_19 <= _GEN_2363;
      end else begin
        REG_7_19 <= _GEN_2395;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_20 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_20 <= _GEN_2524;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_20 <= _GEN_2364;
      end else begin
        REG_7_20 <= _GEN_2396;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_21 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_21 <= _GEN_2525;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_21 <= _GEN_2365;
      end else begin
        REG_7_21 <= _GEN_2397;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_22 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_22 <= _GEN_2526;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_22 <= _GEN_2366;
      end else begin
        REG_7_22 <= _GEN_2398;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_23 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_23 <= _GEN_2527;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_23 <= _GEN_2367;
      end else begin
        REG_7_23 <= _GEN_2399;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_24 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_24 <= _GEN_2528;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_24 <= _GEN_2368;
      end else begin
        REG_7_24 <= _GEN_2400;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_25 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_25 <= _GEN_2529;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_25 <= _GEN_2369;
      end else begin
        REG_7_25 <= _GEN_2401;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_26 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_26 <= _GEN_2530;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_26 <= _GEN_2370;
      end else begin
        REG_7_26 <= _GEN_2402;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_27 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_27 <= _GEN_2531;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_27 <= _GEN_2371;
      end else begin
        REG_7_27 <= _GEN_2403;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_28 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_28 <= _GEN_2532;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_28 <= _GEN_2372;
      end else begin
        REG_7_28 <= _GEN_2404;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_29 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_29 <= _GEN_2533;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_29 <= _GEN_2373;
      end else begin
        REG_7_29 <= _GEN_2405;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_30 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_30 <= _GEN_2534;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_30 <= _GEN_2374;
      end else begin
        REG_7_30 <= _GEN_2406;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 98:44]
      REG_7_31 <= 1'h0; // @[SharedPipelinedCache.scala 98:44]
    end else if (~updateLogic_io_cacheUpdateControl_refill & updateLogic_io_cacheUpdateControl_update & isUpdateWay_7
      ) begin // @[SharedPipelinedCache.scala 123:112]
      REG_7_31 <= _GEN_2535;
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      if (updateLogic_io_cacheUpdateControl_update) begin // @[SharedPipelinedCache.scala 115:54]
        REG_7_31 <= _GEN_2375;
      end else begin
        REG_7_31 <= _GEN_2407;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_0 <= _GEN_72;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_1 <= _GEN_73;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_2 <= _GEN_74;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_3 <= _GEN_75;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_4 <= _GEN_76;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_5 <= _GEN_77;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_6 <= _GEN_78;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_7 <= _GEN_79;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_8 <= _GEN_80;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_9 <= _GEN_81;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_10 <= _GEN_82;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_11 <= _GEN_83;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_12 <= _GEN_84;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_13 <= _GEN_85;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_14 <= _GEN_86;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_15 <= _GEN_87;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_16 <= _GEN_88;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_17 <= _GEN_89;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_18 <= _GEN_90;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_19 <= _GEN_91;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_20 <= _GEN_92;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_21 <= _GEN_93;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_22 <= _GEN_94;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_23 <= _GEN_95;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_24 <= _GEN_96;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_25 <= _GEN_97;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_26 <= _GEN_98;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_27 <= _GEN_99;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_28 <= _GEN_100;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_29 <= _GEN_101;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_30 <= _GEN_102;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_8_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T) begin // @[SharedPipelinedCache.scala 112:67]
      REG_8_31 <= _GEN_103;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_0 <= _GEN_392;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_1 <= _GEN_393;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_2 <= _GEN_394;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_3 <= _GEN_395;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_4 <= _GEN_396;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_5 <= _GEN_397;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_6 <= _GEN_398;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_7 <= _GEN_399;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_8 <= _GEN_400;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_9 <= _GEN_401;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_10 <= _GEN_402;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_11 <= _GEN_403;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_12 <= _GEN_404;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_13 <= _GEN_405;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_14 <= _GEN_406;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_15 <= _GEN_407;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_16 <= _GEN_408;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_17 <= _GEN_409;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_18 <= _GEN_410;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_19 <= _GEN_411;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_20 <= _GEN_412;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_21 <= _GEN_413;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_22 <= _GEN_414;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_23 <= _GEN_415;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_24 <= _GEN_416;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_25 <= _GEN_417;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_26 <= _GEN_418;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_27 <= _GEN_419;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_28 <= _GEN_420;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_29 <= _GEN_421;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_30 <= _GEN_422;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_9_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_1) begin // @[SharedPipelinedCache.scala 112:67]
      REG_9_31 <= _GEN_423;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_0 <= _GEN_712;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_1 <= _GEN_713;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_2 <= _GEN_714;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_3 <= _GEN_715;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_4 <= _GEN_716;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_5 <= _GEN_717;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_6 <= _GEN_718;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_7 <= _GEN_719;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_8 <= _GEN_720;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_9 <= _GEN_721;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_10 <= _GEN_722;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_11 <= _GEN_723;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_12 <= _GEN_724;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_13 <= _GEN_725;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_14 <= _GEN_726;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_15 <= _GEN_727;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_16 <= _GEN_728;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_17 <= _GEN_729;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_18 <= _GEN_730;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_19 <= _GEN_731;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_20 <= _GEN_732;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_21 <= _GEN_733;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_22 <= _GEN_734;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_23 <= _GEN_735;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_24 <= _GEN_736;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_25 <= _GEN_737;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_26 <= _GEN_738;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_27 <= _GEN_739;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_28 <= _GEN_740;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_29 <= _GEN_741;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_30 <= _GEN_742;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_10_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_2) begin // @[SharedPipelinedCache.scala 112:67]
      REG_10_31 <= _GEN_743;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_0 <= _GEN_1032;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_1 <= _GEN_1033;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_2 <= _GEN_1034;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_3 <= _GEN_1035;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_4 <= _GEN_1036;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_5 <= _GEN_1037;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_6 <= _GEN_1038;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_7 <= _GEN_1039;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_8 <= _GEN_1040;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_9 <= _GEN_1041;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_10 <= _GEN_1042;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_11 <= _GEN_1043;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_12 <= _GEN_1044;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_13 <= _GEN_1045;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_14 <= _GEN_1046;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_15 <= _GEN_1047;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_16 <= _GEN_1048;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_17 <= _GEN_1049;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_18 <= _GEN_1050;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_19 <= _GEN_1051;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_20 <= _GEN_1052;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_21 <= _GEN_1053;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_22 <= _GEN_1054;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_23 <= _GEN_1055;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_24 <= _GEN_1056;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_25 <= _GEN_1057;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_26 <= _GEN_1058;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_27 <= _GEN_1059;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_28 <= _GEN_1060;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_29 <= _GEN_1061;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_30 <= _GEN_1062;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_11_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_3) begin // @[SharedPipelinedCache.scala 112:67]
      REG_11_31 <= _GEN_1063;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_0 <= _GEN_1352;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_1 <= _GEN_1353;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_2 <= _GEN_1354;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_3 <= _GEN_1355;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_4 <= _GEN_1356;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_5 <= _GEN_1357;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_6 <= _GEN_1358;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_7 <= _GEN_1359;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_8 <= _GEN_1360;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_9 <= _GEN_1361;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_10 <= _GEN_1362;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_11 <= _GEN_1363;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_12 <= _GEN_1364;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_13 <= _GEN_1365;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_14 <= _GEN_1366;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_15 <= _GEN_1367;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_16 <= _GEN_1368;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_17 <= _GEN_1369;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_18 <= _GEN_1370;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_19 <= _GEN_1371;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_20 <= _GEN_1372;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_21 <= _GEN_1373;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_22 <= _GEN_1374;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_23 <= _GEN_1375;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_24 <= _GEN_1376;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_25 <= _GEN_1377;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_26 <= _GEN_1378;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_27 <= _GEN_1379;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_28 <= _GEN_1380;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_29 <= _GEN_1381;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_30 <= _GEN_1382;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_12_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_4) begin // @[SharedPipelinedCache.scala 112:67]
      REG_12_31 <= _GEN_1383;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_0 <= _GEN_1672;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_1 <= _GEN_1673;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_2 <= _GEN_1674;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_3 <= _GEN_1675;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_4 <= _GEN_1676;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_5 <= _GEN_1677;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_6 <= _GEN_1678;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_7 <= _GEN_1679;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_8 <= _GEN_1680;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_9 <= _GEN_1681;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_10 <= _GEN_1682;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_11 <= _GEN_1683;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_12 <= _GEN_1684;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_13 <= _GEN_1685;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_14 <= _GEN_1686;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_15 <= _GEN_1687;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_16 <= _GEN_1688;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_17 <= _GEN_1689;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_18 <= _GEN_1690;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_19 <= _GEN_1691;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_20 <= _GEN_1692;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_21 <= _GEN_1693;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_22 <= _GEN_1694;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_23 <= _GEN_1695;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_24 <= _GEN_1696;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_25 <= _GEN_1697;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_26 <= _GEN_1698;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_27 <= _GEN_1699;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_28 <= _GEN_1700;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_29 <= _GEN_1701;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_30 <= _GEN_1702;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_13_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_5) begin // @[SharedPipelinedCache.scala 112:67]
      REG_13_31 <= _GEN_1703;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_0 <= _GEN_1992;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_1 <= _GEN_1993;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_2 <= _GEN_1994;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_3 <= _GEN_1995;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_4 <= _GEN_1996;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_5 <= _GEN_1997;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_6 <= _GEN_1998;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_7 <= _GEN_1999;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_8 <= _GEN_2000;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_9 <= _GEN_2001;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_10 <= _GEN_2002;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_11 <= _GEN_2003;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_12 <= _GEN_2004;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_13 <= _GEN_2005;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_14 <= _GEN_2006;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_15 <= _GEN_2007;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_16 <= _GEN_2008;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_17 <= _GEN_2009;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_18 <= _GEN_2010;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_19 <= _GEN_2011;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_20 <= _GEN_2012;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_21 <= _GEN_2013;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_22 <= _GEN_2014;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_23 <= _GEN_2015;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_24 <= _GEN_2016;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_25 <= _GEN_2017;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_26 <= _GEN_2018;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_27 <= _GEN_2019;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_28 <= _GEN_2020;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_29 <= _GEN_2021;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_30 <= _GEN_2022;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_14_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_6) begin // @[SharedPipelinedCache.scala 112:67]
      REG_14_31 <= _GEN_2023;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_0 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_0 <= _GEN_2312;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_1 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_1 <= _GEN_2313;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_2 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_2 <= _GEN_2314;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_3 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_3 <= _GEN_2315;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_4 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_4 <= _GEN_2316;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_5 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_5 <= _GEN_2317;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_6 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_6 <= _GEN_2318;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_7 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_7 <= _GEN_2319;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_8 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_8 <= _GEN_2320;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_9 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_9 <= _GEN_2321;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_10 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_10 <= _GEN_2322;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_11 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_11 <= _GEN_2323;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_12 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_12 <= _GEN_2324;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_13 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_13 <= _GEN_2325;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_14 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_14 <= _GEN_2326;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_15 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_15 <= _GEN_2327;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_16 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_16 <= _GEN_2328;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_17 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_17 <= _GEN_2329;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_18 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_18 <= _GEN_2330;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_19 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_19 <= _GEN_2331;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_20 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_20 <= _GEN_2332;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_21 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_21 <= _GEN_2333;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_22 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_22 <= _GEN_2334;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_23 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_23 <= _GEN_2335;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_24 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_24 <= _GEN_2336;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_25 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_25 <= _GEN_2337;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_26 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_26 <= _GEN_2338;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_27 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_27 <= _GEN_2339;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_28 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_28 <= _GEN_2340;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_29 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_29 <= _GEN_2341;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_30 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_30 <= _GEN_2342;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 99:44]
      REG_15_31 <= 1'h0; // @[SharedPipelinedCache.scala 99:44]
    end else if (_T_7) begin // @[SharedPipelinedCache.scala 112:67]
      REG_15_31 <= _GEN_2343;
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      coreIdRepReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      coreIdRepReg <= coreIdTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqValidRepReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqValidRepReg <= reqValidTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqIdRepReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqIdRepReg <= reqIdTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqRwRepReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqRwRepReg <= reqRwTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      wDataRepReg <= 128'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      wDataRepReg <= wDataTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      hitRepReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      hitRepReg <= hit; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      hitWayRepReg <= 3'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (hits_0) begin // @[Mux.scala 47:70]
        hitWayRepReg <= 3'h0;
      end else if (hits_1) begin // @[Mux.scala 47:70]
        hitWayRepReg <= 3'h1;
      end else begin
        hitWayRepReg <= _hitWay_T_4;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_0 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_0 <= REG__31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_0 <= REG__30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_0 <= _GEN_69;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_1 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_1 <= REG_1_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_1 <= REG_1_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_1 <= _GEN_389;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_2 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_2 <= REG_2_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_2 <= REG_2_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_2 <= _GEN_709;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_3 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_3 <= REG_3_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_3 <= REG_3_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_3 <= _GEN_1029;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_4 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_4 <= REG_4_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_4 <= REG_4_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_4 <= _GEN_1349;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_5 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_5 <= REG_5_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_5 <= REG_5_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_5 <= _GEN_1669;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_6 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_6 <= REG_6_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_6 <= REG_6_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_6 <= _GEN_1989;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyRepReg_7 <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (5'h1f == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_7 <= REG_7_31; // @[SharedPipelinedCache.scala 107:19]
      end else if (5'h1e == indexTagReg) begin // @[SharedPipelinedCache.scala 107:19]
        dirtyRepReg_7 <= REG_7_30; // @[SharedPipelinedCache.scala 107:19]
      end else begin
        dirtyRepReg_7 <= _GEN_2309;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_0 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_0 <= readTags_0; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_1 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_1 <= readTags_1; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_2 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_2 <= readTags_2; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_3 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_3 <= readTags_3; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_4 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_4 <= readTags_4; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_5 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_5 <= readTags_5; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_6 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_6 <= readTags_6; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      readTagsRepReg_7 <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      readTagsRepReg_7 <= readTags_7; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      blockRepReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      blockRepReg <= blockTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      indexRepReg <= 5'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      indexRepReg <= indexTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      tagRepReg <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      tagRepReg <= tagTagReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      coreIdReadReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      coreIdReadReg <= coreIdRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqValidReadReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqValidReadReg <= reqValidRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqIdReadReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqIdReadReg <= reqIdRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      reqRwReadReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      reqRwReadReg <= reqRwRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      wDataReadReg <= 128'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      wDataReadReg <= wDataRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      hitReadReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      hitReadReg <= hitRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      hitWayReadReg <= 3'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      hitWayReadReg <= hitWayRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      isRepDirtyReadReg <= 1'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (3'h7 == io_repPol_replaceWay) begin // @[SharedPipelinedCache.scala 44:19]
        isRepDirtyReadReg <= dirtyRepReg_7; // @[SharedPipelinedCache.scala 44:19]
      end else if (3'h6 == io_repPol_replaceWay) begin // @[SharedPipelinedCache.scala 44:19]
        isRepDirtyReadReg <= dirtyRepReg_6; // @[SharedPipelinedCache.scala 44:19]
      end else begin
        isRepDirtyReadReg <= _GEN_2608;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      dirtyTagReadReg <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      if (3'h7 == io_repPol_replaceWay) begin // @[SharedPipelinedCache.scala 44:19]
        dirtyTagReadReg <= readTagsRepReg_7; // @[SharedPipelinedCache.scala 44:19]
      end else if (3'h6 == io_repPol_replaceWay) begin // @[SharedPipelinedCache.scala 44:19]
        dirtyTagReadReg <= readTagsRepReg_6; // @[SharedPipelinedCache.scala 44:19]
      end else begin
        dirtyTagReadReg <= _GEN_2617;
      end
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      blockReadReg <= 2'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      blockReadReg <= blockRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      indexReadReg <= 5'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      indexReadReg <= indexRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
    if (reset) begin // @[SharedPipelinedCache.scala 42:30]
      tagReadReg <= 4'h0; // @[SharedPipelinedCache.scala 42:30]
    end else if (_reqAccept_T) begin // @[SharedPipelinedCache.scala 43:14]
      tagReadReg <= tagRepReg; // @[SharedPipelinedCache.scala 44:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  coreIdTagReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reqValidTagReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reqIdTagReg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  reqRwTagReg = _RAND_3[0:0];
  _RAND_4 = {4{`RANDOM}};
  wDataTagReg = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  blockTagReg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  indexTagReg = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  tagTagReg = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  REG__0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG__1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG__2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG__3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG__4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG__5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG__6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  REG__7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG__8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG__9 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG__10 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG__11 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG__12 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  REG__13 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  REG__14 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  REG__15 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG__16 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  REG__17 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  REG__18 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG__19 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  REG__20 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  REG__21 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  REG__22 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  REG__23 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  REG__24 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  REG__25 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  REG__26 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  REG__27 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  REG__28 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  REG__29 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  REG__30 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG__31 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG_1_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG_1_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG_1_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG_1_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG_1_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG_1_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_1_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG_1_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG_1_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG_1_9 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG_1_10 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG_1_11 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG_1_12 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  REG_1_13 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  REG_1_14 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  REG_1_15 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  REG_1_16 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  REG_1_17 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  REG_1_18 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  REG_1_19 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  REG_1_20 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  REG_1_21 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  REG_1_22 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  REG_1_23 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  REG_1_24 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  REG_1_25 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  REG_1_26 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  REG_1_27 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  REG_1_28 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  REG_1_29 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  REG_1_30 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  REG_1_31 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  REG_2_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  REG_2_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  REG_2_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  REG_2_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  REG_2_4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  REG_2_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  REG_2_6 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  REG_2_7 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  REG_2_8 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  REG_2_9 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  REG_2_10 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  REG_2_11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  REG_2_12 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  REG_2_13 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  REG_2_14 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  REG_2_15 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  REG_2_16 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  REG_2_17 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG_2_18 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  REG_2_19 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  REG_2_20 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  REG_2_21 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  REG_2_22 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  REG_2_23 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  REG_2_24 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  REG_2_25 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  REG_2_26 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  REG_2_27 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG_2_28 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG_2_29 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  REG_2_30 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  REG_2_31 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG_3_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  REG_3_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  REG_3_2 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG_3_3 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG_3_4 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG_3_5 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  REG_3_6 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  REG_3_7 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG_3_8 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  REG_3_9 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG_3_10 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  REG_3_11 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  REG_3_12 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG_3_13 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG_3_14 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  REG_3_15 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG_3_16 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  REG_3_17 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  REG_3_18 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  REG_3_19 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  REG_3_20 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  REG_3_21 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  REG_3_22 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  REG_3_23 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  REG_3_24 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  REG_3_25 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  REG_3_26 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  REG_3_27 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  REG_3_28 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  REG_3_29 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  REG_3_30 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  REG_3_31 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  REG_4_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  REG_4_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  REG_4_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  REG_4_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  REG_4_4 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  REG_4_5 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  REG_4_6 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  REG_4_7 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  REG_4_8 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  REG_4_9 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  REG_4_10 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  REG_4_11 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  REG_4_12 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  REG_4_13 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  REG_4_14 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  REG_4_15 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  REG_4_16 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  REG_4_17 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  REG_4_18 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  REG_4_19 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  REG_4_20 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  REG_4_21 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  REG_4_22 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  REG_4_23 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  REG_4_24 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  REG_4_25 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  REG_4_26 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  REG_4_27 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  REG_4_28 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  REG_4_29 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  REG_4_30 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  REG_4_31 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  REG_5_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  REG_5_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  REG_5_2 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  REG_5_3 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  REG_5_4 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  REG_5_5 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  REG_5_6 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  REG_5_7 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  REG_5_8 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  REG_5_9 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  REG_5_10 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  REG_5_11 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  REG_5_12 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  REG_5_13 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  REG_5_14 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  REG_5_15 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  REG_5_16 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  REG_5_17 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  REG_5_18 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  REG_5_19 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  REG_5_20 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  REG_5_21 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  REG_5_22 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  REG_5_23 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  REG_5_24 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  REG_5_25 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  REG_5_26 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  REG_5_27 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  REG_5_28 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  REG_5_29 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  REG_5_30 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  REG_5_31 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  REG_6_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  REG_6_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  REG_6_2 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  REG_6_3 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  REG_6_4 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  REG_6_5 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  REG_6_6 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  REG_6_7 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  REG_6_8 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  REG_6_9 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  REG_6_10 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  REG_6_11 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  REG_6_12 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  REG_6_13 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  REG_6_14 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  REG_6_15 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  REG_6_16 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  REG_6_17 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  REG_6_18 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  REG_6_19 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  REG_6_20 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  REG_6_21 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  REG_6_22 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  REG_6_23 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  REG_6_24 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  REG_6_25 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  REG_6_26 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  REG_6_27 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  REG_6_28 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  REG_6_29 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  REG_6_30 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  REG_6_31 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  REG_7_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  REG_7_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  REG_7_2 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  REG_7_3 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  REG_7_4 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  REG_7_5 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  REG_7_6 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  REG_7_7 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  REG_7_8 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  REG_7_9 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  REG_7_10 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  REG_7_11 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  REG_7_12 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  REG_7_13 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  REG_7_14 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  REG_7_15 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  REG_7_16 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  REG_7_17 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  REG_7_18 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  REG_7_19 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  REG_7_20 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  REG_7_21 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  REG_7_22 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  REG_7_23 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  REG_7_24 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  REG_7_25 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  REG_7_26 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  REG_7_27 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  REG_7_28 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  REG_7_29 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  REG_7_30 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  REG_7_31 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  REG_8_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  REG_8_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  REG_8_2 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  REG_8_3 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  REG_8_4 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  REG_8_5 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  REG_8_6 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  REG_8_7 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  REG_8_8 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  REG_8_9 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  REG_8_10 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  REG_8_11 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  REG_8_12 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  REG_8_13 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  REG_8_14 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  REG_8_15 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  REG_8_16 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  REG_8_17 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  REG_8_18 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  REG_8_19 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  REG_8_20 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  REG_8_21 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  REG_8_22 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  REG_8_23 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  REG_8_24 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  REG_8_25 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  REG_8_26 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  REG_8_27 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  REG_8_28 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  REG_8_29 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  REG_8_30 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  REG_8_31 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  REG_9_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  REG_9_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  REG_9_2 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  REG_9_3 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  REG_9_4 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  REG_9_5 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  REG_9_6 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  REG_9_7 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  REG_9_8 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  REG_9_9 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  REG_9_10 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  REG_9_11 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  REG_9_12 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  REG_9_13 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  REG_9_14 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  REG_9_15 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  REG_9_16 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  REG_9_17 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  REG_9_18 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  REG_9_19 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  REG_9_20 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  REG_9_21 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  REG_9_22 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  REG_9_23 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  REG_9_24 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  REG_9_25 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  REG_9_26 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  REG_9_27 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  REG_9_28 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  REG_9_29 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  REG_9_30 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  REG_9_31 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  REG_10_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  REG_10_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  REG_10_2 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  REG_10_3 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  REG_10_4 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  REG_10_5 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  REG_10_6 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  REG_10_7 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  REG_10_8 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  REG_10_9 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  REG_10_10 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  REG_10_11 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  REG_10_12 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  REG_10_13 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  REG_10_14 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  REG_10_15 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  REG_10_16 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  REG_10_17 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  REG_10_18 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  REG_10_19 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  REG_10_20 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  REG_10_21 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  REG_10_22 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  REG_10_23 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  REG_10_24 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  REG_10_25 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  REG_10_26 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  REG_10_27 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  REG_10_28 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  REG_10_29 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  REG_10_30 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  REG_10_31 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  REG_11_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  REG_11_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  REG_11_2 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  REG_11_3 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  REG_11_4 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  REG_11_5 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  REG_11_6 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  REG_11_7 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  REG_11_8 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  REG_11_9 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  REG_11_10 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  REG_11_11 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  REG_11_12 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  REG_11_13 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  REG_11_14 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  REG_11_15 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  REG_11_16 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  REG_11_17 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  REG_11_18 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  REG_11_19 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  REG_11_20 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  REG_11_21 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  REG_11_22 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  REG_11_23 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  REG_11_24 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  REG_11_25 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  REG_11_26 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  REG_11_27 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  REG_11_28 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  REG_11_29 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  REG_11_30 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  REG_11_31 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  REG_12_0 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  REG_12_1 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  REG_12_2 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  REG_12_3 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  REG_12_4 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  REG_12_5 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  REG_12_6 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  REG_12_7 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  REG_12_8 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  REG_12_9 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  REG_12_10 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  REG_12_11 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  REG_12_12 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  REG_12_13 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  REG_12_14 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  REG_12_15 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  REG_12_16 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  REG_12_17 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  REG_12_18 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  REG_12_19 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  REG_12_20 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  REG_12_21 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  REG_12_22 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  REG_12_23 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  REG_12_24 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  REG_12_25 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  REG_12_26 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  REG_12_27 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  REG_12_28 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  REG_12_29 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  REG_12_30 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  REG_12_31 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  REG_13_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  REG_13_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  REG_13_2 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  REG_13_3 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  REG_13_4 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  REG_13_5 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  REG_13_6 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  REG_13_7 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  REG_13_8 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  REG_13_9 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  REG_13_10 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  REG_13_11 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  REG_13_12 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  REG_13_13 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  REG_13_14 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  REG_13_15 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  REG_13_16 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  REG_13_17 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  REG_13_18 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  REG_13_19 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  REG_13_20 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  REG_13_21 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  REG_13_22 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  REG_13_23 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  REG_13_24 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  REG_13_25 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  REG_13_26 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  REG_13_27 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  REG_13_28 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  REG_13_29 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  REG_13_30 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  REG_13_31 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  REG_14_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  REG_14_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  REG_14_2 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  REG_14_3 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  REG_14_4 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  REG_14_5 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  REG_14_6 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  REG_14_7 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  REG_14_8 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  REG_14_9 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  REG_14_10 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  REG_14_11 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  REG_14_12 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  REG_14_13 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  REG_14_14 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  REG_14_15 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  REG_14_16 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  REG_14_17 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  REG_14_18 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  REG_14_19 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  REG_14_20 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  REG_14_21 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  REG_14_22 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  REG_14_23 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  REG_14_24 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  REG_14_25 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  REG_14_26 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  REG_14_27 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  REG_14_28 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  REG_14_29 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  REG_14_30 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  REG_14_31 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  REG_15_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  REG_15_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  REG_15_2 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  REG_15_3 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  REG_15_4 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  REG_15_5 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  REG_15_6 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  REG_15_7 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  REG_15_8 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  REG_15_9 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  REG_15_10 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  REG_15_11 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  REG_15_12 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  REG_15_13 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  REG_15_14 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  REG_15_15 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  REG_15_16 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  REG_15_17 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  REG_15_18 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  REG_15_19 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  REG_15_20 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  REG_15_21 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  REG_15_22 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  REG_15_23 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  REG_15_24 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  REG_15_25 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  REG_15_26 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  REG_15_27 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  REG_15_28 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  REG_15_29 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  REG_15_30 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  REG_15_31 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  coreIdRepReg = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  reqValidRepReg = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  reqIdRepReg = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  reqRwRepReg = _RAND_523[0:0];
  _RAND_524 = {4{`RANDOM}};
  wDataRepReg = _RAND_524[127:0];
  _RAND_525 = {1{`RANDOM}};
  hitRepReg = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  hitWayRepReg = _RAND_526[2:0];
  _RAND_527 = {1{`RANDOM}};
  dirtyRepReg_0 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  dirtyRepReg_1 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  dirtyRepReg_2 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dirtyRepReg_3 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  dirtyRepReg_4 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  dirtyRepReg_5 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dirtyRepReg_6 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  dirtyRepReg_7 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  readTagsRepReg_0 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  readTagsRepReg_1 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  readTagsRepReg_2 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  readTagsRepReg_3 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  readTagsRepReg_4 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  readTagsRepReg_5 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  readTagsRepReg_6 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  readTagsRepReg_7 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  blockRepReg = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  indexRepReg = _RAND_544[4:0];
  _RAND_545 = {1{`RANDOM}};
  tagRepReg = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  coreIdReadReg = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  reqValidReadReg = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  reqIdReadReg = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  reqRwReadReg = _RAND_549[0:0];
  _RAND_550 = {4{`RANDOM}};
  wDataReadReg = _RAND_550[127:0];
  _RAND_551 = {1{`RANDOM}};
  hitReadReg = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  hitWayReadReg = _RAND_552[2:0];
  _RAND_553 = {1{`RANDOM}};
  isRepDirtyReadReg = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dirtyTagReadReg = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  blockReadReg = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  indexReadReg = _RAND_556[4:0];
  _RAND_557 = {1{`RANDOM}};
  tagReadReg = _RAND_557[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BitPlruReplacementPolicy(
  input        clock,
  input        reset,
  input        io_control_update_valid,
  input  [2:0] io_control_update_bits,
  input        io_control_stall,
  input  [4:0] io_control_setIdx,
  output [2:0] io_control_replaceWay
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
`endif // RANDOMIZE_REG_INIT
  reg  REG__0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG__7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_1_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_2_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_3_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_4_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_5_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_6_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_7_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_8_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_9_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_10_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_11_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_12_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_13_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_14_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_15_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_16_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_17_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_18_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_19_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_20_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_21_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_22_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_23_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_24_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_25_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_26_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_27_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_28_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_29_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_30_7; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_0; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_1; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_2; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_3; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_4; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_5; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_6; // @[BitPlruReplacementPolicy.scala 87:45]
  reg  REG_31_7; // @[BitPlruReplacementPolicy.scala 87:45]
  wire  _GEN_15 = 5'h0 == io_control_setIdx & REG__7; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_39 = 5'h1 == io_control_setIdx ? REG_1_7 : _GEN_15; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_63 = 5'h2 == io_control_setIdx ? REG_2_7 : _GEN_39; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_87 = 5'h3 == io_control_setIdx ? REG_3_7 : _GEN_63; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_111 = 5'h4 == io_control_setIdx ? REG_4_7 : _GEN_87; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_135 = 5'h5 == io_control_setIdx ? REG_5_7 : _GEN_111; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_159 = 5'h6 == io_control_setIdx ? REG_6_7 : _GEN_135; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_183 = 5'h7 == io_control_setIdx ? REG_7_7 : _GEN_159; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_207 = 5'h8 == io_control_setIdx ? REG_8_7 : _GEN_183; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_231 = 5'h9 == io_control_setIdx ? REG_9_7 : _GEN_207; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_255 = 5'ha == io_control_setIdx ? REG_10_7 : _GEN_231; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_279 = 5'hb == io_control_setIdx ? REG_11_7 : _GEN_255; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_303 = 5'hc == io_control_setIdx ? REG_12_7 : _GEN_279; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_327 = 5'hd == io_control_setIdx ? REG_13_7 : _GEN_303; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_351 = 5'he == io_control_setIdx ? REG_14_7 : _GEN_327; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_375 = 5'hf == io_control_setIdx ? REG_15_7 : _GEN_351; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_399 = 5'h10 == io_control_setIdx ? REG_16_7 : _GEN_375; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_423 = 5'h11 == io_control_setIdx ? REG_17_7 : _GEN_399; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_447 = 5'h12 == io_control_setIdx ? REG_18_7 : _GEN_423; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_471 = 5'h13 == io_control_setIdx ? REG_19_7 : _GEN_447; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_495 = 5'h14 == io_control_setIdx ? REG_20_7 : _GEN_471; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_519 = 5'h15 == io_control_setIdx ? REG_21_7 : _GEN_495; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_543 = 5'h16 == io_control_setIdx ? REG_22_7 : _GEN_519; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_567 = 5'h17 == io_control_setIdx ? REG_23_7 : _GEN_543; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_591 = 5'h18 == io_control_setIdx ? REG_24_7 : _GEN_567; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_615 = 5'h19 == io_control_setIdx ? REG_25_7 : _GEN_591; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_639 = 5'h1a == io_control_setIdx ? REG_26_7 : _GEN_615; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_663 = 5'h1b == io_control_setIdx ? REG_27_7 : _GEN_639; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_687 = 5'h1c == io_control_setIdx ? REG_28_7 : _GEN_663; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_711 = 5'h1d == io_control_setIdx ? REG_29_7 : _GEN_687; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_735 = 5'h1e == io_control_setIdx ? REG_30_7 : _GEN_711; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_7 = 5'h1f == io_control_setIdx ? REG_31_7 : _GEN_735; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_14 = 5'h0 == io_control_setIdx & REG__6; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_38 = 5'h1 == io_control_setIdx ? REG_1_6 : _GEN_14; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_62 = 5'h2 == io_control_setIdx ? REG_2_6 : _GEN_38; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_86 = 5'h3 == io_control_setIdx ? REG_3_6 : _GEN_62; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_110 = 5'h4 == io_control_setIdx ? REG_4_6 : _GEN_86; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_134 = 5'h5 == io_control_setIdx ? REG_5_6 : _GEN_110; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_158 = 5'h6 == io_control_setIdx ? REG_6_6 : _GEN_134; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_182 = 5'h7 == io_control_setIdx ? REG_7_6 : _GEN_158; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_206 = 5'h8 == io_control_setIdx ? REG_8_6 : _GEN_182; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_230 = 5'h9 == io_control_setIdx ? REG_9_6 : _GEN_206; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_254 = 5'ha == io_control_setIdx ? REG_10_6 : _GEN_230; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_278 = 5'hb == io_control_setIdx ? REG_11_6 : _GEN_254; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_302 = 5'hc == io_control_setIdx ? REG_12_6 : _GEN_278; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_326 = 5'hd == io_control_setIdx ? REG_13_6 : _GEN_302; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_350 = 5'he == io_control_setIdx ? REG_14_6 : _GEN_326; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_374 = 5'hf == io_control_setIdx ? REG_15_6 : _GEN_350; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_398 = 5'h10 == io_control_setIdx ? REG_16_6 : _GEN_374; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_422 = 5'h11 == io_control_setIdx ? REG_17_6 : _GEN_398; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_446 = 5'h12 == io_control_setIdx ? REG_18_6 : _GEN_422; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_470 = 5'h13 == io_control_setIdx ? REG_19_6 : _GEN_446; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_494 = 5'h14 == io_control_setIdx ? REG_20_6 : _GEN_470; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_518 = 5'h15 == io_control_setIdx ? REG_21_6 : _GEN_494; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_542 = 5'h16 == io_control_setIdx ? REG_22_6 : _GEN_518; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_566 = 5'h17 == io_control_setIdx ? REG_23_6 : _GEN_542; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_590 = 5'h18 == io_control_setIdx ? REG_24_6 : _GEN_566; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_614 = 5'h19 == io_control_setIdx ? REG_25_6 : _GEN_590; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_638 = 5'h1a == io_control_setIdx ? REG_26_6 : _GEN_614; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_662 = 5'h1b == io_control_setIdx ? REG_27_6 : _GEN_638; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_686 = 5'h1c == io_control_setIdx ? REG_28_6 : _GEN_662; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_710 = 5'h1d == io_control_setIdx ? REG_29_6 : _GEN_686; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_734 = 5'h1e == io_control_setIdx ? REG_30_6 : _GEN_710; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_6 = 5'h1f == io_control_setIdx ? REG_31_6 : _GEN_734; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_13 = 5'h0 == io_control_setIdx & REG__5; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_37 = 5'h1 == io_control_setIdx ? REG_1_5 : _GEN_13; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_61 = 5'h2 == io_control_setIdx ? REG_2_5 : _GEN_37; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_85 = 5'h3 == io_control_setIdx ? REG_3_5 : _GEN_61; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_109 = 5'h4 == io_control_setIdx ? REG_4_5 : _GEN_85; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_133 = 5'h5 == io_control_setIdx ? REG_5_5 : _GEN_109; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_157 = 5'h6 == io_control_setIdx ? REG_6_5 : _GEN_133; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_181 = 5'h7 == io_control_setIdx ? REG_7_5 : _GEN_157; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_205 = 5'h8 == io_control_setIdx ? REG_8_5 : _GEN_181; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_229 = 5'h9 == io_control_setIdx ? REG_9_5 : _GEN_205; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_253 = 5'ha == io_control_setIdx ? REG_10_5 : _GEN_229; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_277 = 5'hb == io_control_setIdx ? REG_11_5 : _GEN_253; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_301 = 5'hc == io_control_setIdx ? REG_12_5 : _GEN_277; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_325 = 5'hd == io_control_setIdx ? REG_13_5 : _GEN_301; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_349 = 5'he == io_control_setIdx ? REG_14_5 : _GEN_325; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_373 = 5'hf == io_control_setIdx ? REG_15_5 : _GEN_349; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_397 = 5'h10 == io_control_setIdx ? REG_16_5 : _GEN_373; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_421 = 5'h11 == io_control_setIdx ? REG_17_5 : _GEN_397; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_445 = 5'h12 == io_control_setIdx ? REG_18_5 : _GEN_421; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_469 = 5'h13 == io_control_setIdx ? REG_19_5 : _GEN_445; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_493 = 5'h14 == io_control_setIdx ? REG_20_5 : _GEN_469; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_517 = 5'h15 == io_control_setIdx ? REG_21_5 : _GEN_493; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_541 = 5'h16 == io_control_setIdx ? REG_22_5 : _GEN_517; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_565 = 5'h17 == io_control_setIdx ? REG_23_5 : _GEN_541; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_589 = 5'h18 == io_control_setIdx ? REG_24_5 : _GEN_565; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_613 = 5'h19 == io_control_setIdx ? REG_25_5 : _GEN_589; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_637 = 5'h1a == io_control_setIdx ? REG_26_5 : _GEN_613; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_661 = 5'h1b == io_control_setIdx ? REG_27_5 : _GEN_637; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_685 = 5'h1c == io_control_setIdx ? REG_28_5 : _GEN_661; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_709 = 5'h1d == io_control_setIdx ? REG_29_5 : _GEN_685; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_733 = 5'h1e == io_control_setIdx ? REG_30_5 : _GEN_709; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_5 = 5'h1f == io_control_setIdx ? REG_31_5 : _GEN_733; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_12 = 5'h0 == io_control_setIdx & REG__4; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_36 = 5'h1 == io_control_setIdx ? REG_1_4 : _GEN_12; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_60 = 5'h2 == io_control_setIdx ? REG_2_4 : _GEN_36; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_84 = 5'h3 == io_control_setIdx ? REG_3_4 : _GEN_60; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_108 = 5'h4 == io_control_setIdx ? REG_4_4 : _GEN_84; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_132 = 5'h5 == io_control_setIdx ? REG_5_4 : _GEN_108; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_156 = 5'h6 == io_control_setIdx ? REG_6_4 : _GEN_132; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_180 = 5'h7 == io_control_setIdx ? REG_7_4 : _GEN_156; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_204 = 5'h8 == io_control_setIdx ? REG_8_4 : _GEN_180; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_228 = 5'h9 == io_control_setIdx ? REG_9_4 : _GEN_204; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_252 = 5'ha == io_control_setIdx ? REG_10_4 : _GEN_228; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_276 = 5'hb == io_control_setIdx ? REG_11_4 : _GEN_252; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_300 = 5'hc == io_control_setIdx ? REG_12_4 : _GEN_276; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_324 = 5'hd == io_control_setIdx ? REG_13_4 : _GEN_300; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_348 = 5'he == io_control_setIdx ? REG_14_4 : _GEN_324; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_372 = 5'hf == io_control_setIdx ? REG_15_4 : _GEN_348; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_396 = 5'h10 == io_control_setIdx ? REG_16_4 : _GEN_372; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_420 = 5'h11 == io_control_setIdx ? REG_17_4 : _GEN_396; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_444 = 5'h12 == io_control_setIdx ? REG_18_4 : _GEN_420; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_468 = 5'h13 == io_control_setIdx ? REG_19_4 : _GEN_444; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_492 = 5'h14 == io_control_setIdx ? REG_20_4 : _GEN_468; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_516 = 5'h15 == io_control_setIdx ? REG_21_4 : _GEN_492; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_540 = 5'h16 == io_control_setIdx ? REG_22_4 : _GEN_516; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_564 = 5'h17 == io_control_setIdx ? REG_23_4 : _GEN_540; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_588 = 5'h18 == io_control_setIdx ? REG_24_4 : _GEN_564; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_612 = 5'h19 == io_control_setIdx ? REG_25_4 : _GEN_588; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_636 = 5'h1a == io_control_setIdx ? REG_26_4 : _GEN_612; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_660 = 5'h1b == io_control_setIdx ? REG_27_4 : _GEN_636; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_684 = 5'h1c == io_control_setIdx ? REG_28_4 : _GEN_660; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_708 = 5'h1d == io_control_setIdx ? REG_29_4 : _GEN_684; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_732 = 5'h1e == io_control_setIdx ? REG_30_4 : _GEN_708; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_4 = 5'h1f == io_control_setIdx ? REG_31_4 : _GEN_732; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_11 = 5'h0 == io_control_setIdx & REG__3; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_35 = 5'h1 == io_control_setIdx ? REG_1_3 : _GEN_11; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_59 = 5'h2 == io_control_setIdx ? REG_2_3 : _GEN_35; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_83 = 5'h3 == io_control_setIdx ? REG_3_3 : _GEN_59; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_107 = 5'h4 == io_control_setIdx ? REG_4_3 : _GEN_83; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_131 = 5'h5 == io_control_setIdx ? REG_5_3 : _GEN_107; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_155 = 5'h6 == io_control_setIdx ? REG_6_3 : _GEN_131; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_179 = 5'h7 == io_control_setIdx ? REG_7_3 : _GEN_155; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_203 = 5'h8 == io_control_setIdx ? REG_8_3 : _GEN_179; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_227 = 5'h9 == io_control_setIdx ? REG_9_3 : _GEN_203; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_251 = 5'ha == io_control_setIdx ? REG_10_3 : _GEN_227; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_275 = 5'hb == io_control_setIdx ? REG_11_3 : _GEN_251; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_299 = 5'hc == io_control_setIdx ? REG_12_3 : _GEN_275; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_323 = 5'hd == io_control_setIdx ? REG_13_3 : _GEN_299; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_347 = 5'he == io_control_setIdx ? REG_14_3 : _GEN_323; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_371 = 5'hf == io_control_setIdx ? REG_15_3 : _GEN_347; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_395 = 5'h10 == io_control_setIdx ? REG_16_3 : _GEN_371; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_419 = 5'h11 == io_control_setIdx ? REG_17_3 : _GEN_395; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_443 = 5'h12 == io_control_setIdx ? REG_18_3 : _GEN_419; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_467 = 5'h13 == io_control_setIdx ? REG_19_3 : _GEN_443; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_491 = 5'h14 == io_control_setIdx ? REG_20_3 : _GEN_467; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_515 = 5'h15 == io_control_setIdx ? REG_21_3 : _GEN_491; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_539 = 5'h16 == io_control_setIdx ? REG_22_3 : _GEN_515; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_563 = 5'h17 == io_control_setIdx ? REG_23_3 : _GEN_539; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_587 = 5'h18 == io_control_setIdx ? REG_24_3 : _GEN_563; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_611 = 5'h19 == io_control_setIdx ? REG_25_3 : _GEN_587; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_635 = 5'h1a == io_control_setIdx ? REG_26_3 : _GEN_611; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_659 = 5'h1b == io_control_setIdx ? REG_27_3 : _GEN_635; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_683 = 5'h1c == io_control_setIdx ? REG_28_3 : _GEN_659; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_707 = 5'h1d == io_control_setIdx ? REG_29_3 : _GEN_683; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_731 = 5'h1e == io_control_setIdx ? REG_30_3 : _GEN_707; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_3 = 5'h1f == io_control_setIdx ? REG_31_3 : _GEN_731; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_10 = 5'h0 == io_control_setIdx & REG__2; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_34 = 5'h1 == io_control_setIdx ? REG_1_2 : _GEN_10; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_58 = 5'h2 == io_control_setIdx ? REG_2_2 : _GEN_34; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_82 = 5'h3 == io_control_setIdx ? REG_3_2 : _GEN_58; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_106 = 5'h4 == io_control_setIdx ? REG_4_2 : _GEN_82; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_130 = 5'h5 == io_control_setIdx ? REG_5_2 : _GEN_106; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_154 = 5'h6 == io_control_setIdx ? REG_6_2 : _GEN_130; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_178 = 5'h7 == io_control_setIdx ? REG_7_2 : _GEN_154; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_202 = 5'h8 == io_control_setIdx ? REG_8_2 : _GEN_178; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_226 = 5'h9 == io_control_setIdx ? REG_9_2 : _GEN_202; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_250 = 5'ha == io_control_setIdx ? REG_10_2 : _GEN_226; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_274 = 5'hb == io_control_setIdx ? REG_11_2 : _GEN_250; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_298 = 5'hc == io_control_setIdx ? REG_12_2 : _GEN_274; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_322 = 5'hd == io_control_setIdx ? REG_13_2 : _GEN_298; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_346 = 5'he == io_control_setIdx ? REG_14_2 : _GEN_322; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_370 = 5'hf == io_control_setIdx ? REG_15_2 : _GEN_346; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_394 = 5'h10 == io_control_setIdx ? REG_16_2 : _GEN_370; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_418 = 5'h11 == io_control_setIdx ? REG_17_2 : _GEN_394; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_442 = 5'h12 == io_control_setIdx ? REG_18_2 : _GEN_418; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_466 = 5'h13 == io_control_setIdx ? REG_19_2 : _GEN_442; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_490 = 5'h14 == io_control_setIdx ? REG_20_2 : _GEN_466; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_514 = 5'h15 == io_control_setIdx ? REG_21_2 : _GEN_490; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_538 = 5'h16 == io_control_setIdx ? REG_22_2 : _GEN_514; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_562 = 5'h17 == io_control_setIdx ? REG_23_2 : _GEN_538; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_586 = 5'h18 == io_control_setIdx ? REG_24_2 : _GEN_562; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_610 = 5'h19 == io_control_setIdx ? REG_25_2 : _GEN_586; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_634 = 5'h1a == io_control_setIdx ? REG_26_2 : _GEN_610; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_658 = 5'h1b == io_control_setIdx ? REG_27_2 : _GEN_634; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_682 = 5'h1c == io_control_setIdx ? REG_28_2 : _GEN_658; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_706 = 5'h1d == io_control_setIdx ? REG_29_2 : _GEN_682; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_730 = 5'h1e == io_control_setIdx ? REG_30_2 : _GEN_706; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_2 = 5'h1f == io_control_setIdx ? REG_31_2 : _GEN_730; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_9 = 5'h0 == io_control_setIdx & REG__1; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_33 = 5'h1 == io_control_setIdx ? REG_1_1 : _GEN_9; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_57 = 5'h2 == io_control_setIdx ? REG_2_1 : _GEN_33; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_81 = 5'h3 == io_control_setIdx ? REG_3_1 : _GEN_57; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_105 = 5'h4 == io_control_setIdx ? REG_4_1 : _GEN_81; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_129 = 5'h5 == io_control_setIdx ? REG_5_1 : _GEN_105; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_153 = 5'h6 == io_control_setIdx ? REG_6_1 : _GEN_129; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_177 = 5'h7 == io_control_setIdx ? REG_7_1 : _GEN_153; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_201 = 5'h8 == io_control_setIdx ? REG_8_1 : _GEN_177; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_225 = 5'h9 == io_control_setIdx ? REG_9_1 : _GEN_201; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_249 = 5'ha == io_control_setIdx ? REG_10_1 : _GEN_225; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_273 = 5'hb == io_control_setIdx ? REG_11_1 : _GEN_249; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_297 = 5'hc == io_control_setIdx ? REG_12_1 : _GEN_273; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_321 = 5'hd == io_control_setIdx ? REG_13_1 : _GEN_297; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_345 = 5'he == io_control_setIdx ? REG_14_1 : _GEN_321; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_369 = 5'hf == io_control_setIdx ? REG_15_1 : _GEN_345; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_393 = 5'h10 == io_control_setIdx ? REG_16_1 : _GEN_369; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_417 = 5'h11 == io_control_setIdx ? REG_17_1 : _GEN_393; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_441 = 5'h12 == io_control_setIdx ? REG_18_1 : _GEN_417; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_465 = 5'h13 == io_control_setIdx ? REG_19_1 : _GEN_441; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_489 = 5'h14 == io_control_setIdx ? REG_20_1 : _GEN_465; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_513 = 5'h15 == io_control_setIdx ? REG_21_1 : _GEN_489; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_537 = 5'h16 == io_control_setIdx ? REG_22_1 : _GEN_513; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_561 = 5'h17 == io_control_setIdx ? REG_23_1 : _GEN_537; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_585 = 5'h18 == io_control_setIdx ? REG_24_1 : _GEN_561; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_609 = 5'h19 == io_control_setIdx ? REG_25_1 : _GEN_585; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_633 = 5'h1a == io_control_setIdx ? REG_26_1 : _GEN_609; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_657 = 5'h1b == io_control_setIdx ? REG_27_1 : _GEN_633; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_681 = 5'h1c == io_control_setIdx ? REG_28_1 : _GEN_657; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_705 = 5'h1d == io_control_setIdx ? REG_29_1 : _GEN_681; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_729 = 5'h1e == io_control_setIdx ? REG_30_1 : _GEN_705; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_1 = 5'h1f == io_control_setIdx ? REG_31_1 : _GEN_729; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_8 = 5'h0 == io_control_setIdx & REG__0; // @[BitPlruReplacementPolicy.scala 93:41 94:18 89:27]
  wire  _GEN_32 = 5'h1 == io_control_setIdx ? REG_1_0 : _GEN_8; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_56 = 5'h2 == io_control_setIdx ? REG_2_0 : _GEN_32; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_80 = 5'h3 == io_control_setIdx ? REG_3_0 : _GEN_56; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_104 = 5'h4 == io_control_setIdx ? REG_4_0 : _GEN_80; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_128 = 5'h5 == io_control_setIdx ? REG_5_0 : _GEN_104; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_152 = 5'h6 == io_control_setIdx ? REG_6_0 : _GEN_128; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_176 = 5'h7 == io_control_setIdx ? REG_7_0 : _GEN_152; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_200 = 5'h8 == io_control_setIdx ? REG_8_0 : _GEN_176; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_224 = 5'h9 == io_control_setIdx ? REG_9_0 : _GEN_200; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_248 = 5'ha == io_control_setIdx ? REG_10_0 : _GEN_224; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_272 = 5'hb == io_control_setIdx ? REG_11_0 : _GEN_248; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_296 = 5'hc == io_control_setIdx ? REG_12_0 : _GEN_272; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_320 = 5'hd == io_control_setIdx ? REG_13_0 : _GEN_296; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_344 = 5'he == io_control_setIdx ? REG_14_0 : _GEN_320; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_368 = 5'hf == io_control_setIdx ? REG_15_0 : _GEN_344; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_392 = 5'h10 == io_control_setIdx ? REG_16_0 : _GEN_368; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_416 = 5'h11 == io_control_setIdx ? REG_17_0 : _GEN_392; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_440 = 5'h12 == io_control_setIdx ? REG_18_0 : _GEN_416; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_464 = 5'h13 == io_control_setIdx ? REG_19_0 : _GEN_440; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_488 = 5'h14 == io_control_setIdx ? REG_20_0 : _GEN_464; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_512 = 5'h15 == io_control_setIdx ? REG_21_0 : _GEN_488; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_536 = 5'h16 == io_control_setIdx ? REG_22_0 : _GEN_512; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_560 = 5'h17 == io_control_setIdx ? REG_23_0 : _GEN_536; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_584 = 5'h18 == io_control_setIdx ? REG_24_0 : _GEN_560; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_608 = 5'h19 == io_control_setIdx ? REG_25_0 : _GEN_584; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_632 = 5'h1a == io_control_setIdx ? REG_26_0 : _GEN_608; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_656 = 5'h1b == io_control_setIdx ? REG_27_0 : _GEN_632; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_680 = 5'h1c == io_control_setIdx ? REG_28_0 : _GEN_656; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_704 = 5'h1d == io_control_setIdx ? REG_29_0 : _GEN_680; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  _GEN_728 = 5'h1e == io_control_setIdx ? REG_30_0 : _GEN_704; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire  selMruBits_0 = 5'h1f == io_control_setIdx ? REG_31_0 : _GEN_728; // @[BitPlruReplacementPolicy.scala 93:41 94:18]
  wire [7:0] _capacity_T = {selMruBits_7,selMruBits_6,selMruBits_5,selMruBits_4,selMruBits_3,selMruBits_2,selMruBits_1,
    selMruBits_0}; // @[BitPlruReplacementPolicy.scala 21:38]
  wire [7:0] _capacity_T_1 = ~_capacity_T; // @[BitPlruReplacementPolicy.scala 21:22]
  wire [7:0] _capacity_T_5 = _capacity_T_1 - 8'h1; // @[BitPlruReplacementPolicy.scala 21:88]
  wire [7:0] _capacity_T_6 = _capacity_T_1 & _capacity_T_5; // @[BitPlruReplacementPolicy.scala 21:53]
  wire  capacity = _capacity_T_6 == 8'h0; // @[BitPlruReplacementPolicy.scala 21:96]
  wire  _GEN_768 = capacity & 3'h0 != io_control_update_bits ? ~selMruBits_0 : selMruBits_0; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_0 = 3'h0 == io_control_update_bits | _GEN_768; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_769 = capacity & 3'h1 != io_control_update_bits ? ~selMruBits_1 : selMruBits_1; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_1 = 3'h1 == io_control_update_bits | _GEN_769; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_770 = capacity & 3'h2 != io_control_update_bits ? ~selMruBits_2 : selMruBits_2; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_2 = 3'h2 == io_control_update_bits | _GEN_770; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_771 = capacity & 3'h3 != io_control_update_bits ? ~selMruBits_3 : selMruBits_3; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_3 = 3'h3 == io_control_update_bits | _GEN_771; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_772 = capacity & 3'h4 != io_control_update_bits ? ~selMruBits_4 : selMruBits_4; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_4 = 3'h4 == io_control_update_bits | _GEN_772; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_773 = capacity & 3'h5 != io_control_update_bits ? ~selMruBits_5 : selMruBits_5; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_5 = 3'h5 == io_control_update_bits | _GEN_773; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_774 = capacity & 3'h6 != io_control_update_bits ? ~selMruBits_6 : selMruBits_6; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_6 = 3'h6 == io_control_update_bits | _GEN_774; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire  _GEN_775 = capacity & 3'h7 != io_control_update_bits ? ~selMruBits_7 : selMruBits_7; // @[BitPlruReplacementPolicy.scala 24:51 25:28 27:28]
  wire  newMruBits_7 = 3'h7 == io_control_update_bits | _GEN_775; // @[BitPlruReplacementPolicy.scala 31:{21,21}]
  wire [2:0] _replaceWay_T_10 = _capacity_T_1[6] ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _replaceWay_T_11 = _capacity_T_1[5] ? 3'h5 : _replaceWay_T_10; // @[Mux.scala 47:70]
  wire [2:0] _replaceWay_T_12 = _capacity_T_1[4] ? 3'h4 : _replaceWay_T_11; // @[Mux.scala 47:70]
  wire [2:0] _replaceWay_T_13 = _capacity_T_1[3] ? 3'h3 : _replaceWay_T_12; // @[Mux.scala 47:70]
  wire [2:0] _replaceWay_T_14 = _capacity_T_1[2] ? 3'h2 : _replaceWay_T_13; // @[Mux.scala 47:70]
  wire  _replaceWayPipeReg_T = ~io_control_stall; // @[BitPlruReplacementPolicy.scala 109:56]
  reg [2:0] replaceWayPipeReg; // @[SharedCacheReplacementPolicyType.scala 40:30]
  assign io_control_replaceWay = replaceWayPipeReg; // @[BitPlruReplacementPolicy.scala 112:25]
  always @(posedge clock) begin
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG__7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h0 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG__7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_1_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_1_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_2_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h2 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_2_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_3_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h3 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_3_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_4_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h4 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_4_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_5_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h5 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_5_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_6_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h6 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_6_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_7_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h7 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_7_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_8_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h8 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_8_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_9_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h9 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_9_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_10_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'ha == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_10_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_11_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hb == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_11_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_12_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hc == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_12_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_13_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hd == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_13_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_14_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'he == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_14_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_15_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'hf == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_15_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_16_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h10 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_16_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_17_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h11 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_17_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_18_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h12 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_18_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_19_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h13 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_19_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_20_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h14 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_20_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_21_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h15 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_21_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_22_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h16 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_22_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_23_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h17 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_23_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_24_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h18 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_24_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_25_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h19 == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_25_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_26_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1a == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_26_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_27_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1b == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_27_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_28_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1c == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_28_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_29_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1d == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_29_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_30_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1e == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_30_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_0 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_0 <= newMruBits_0; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_1 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_1 <= newMruBits_1; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_2 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_2 <= newMruBits_2; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_3 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_3 <= newMruBits_3; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_4 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_4 <= newMruBits_4; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_5 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_5 <= newMruBits_5; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_6 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_6 <= newMruBits_6; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[BitPlruReplacementPolicy.scala 87:45]
      REG_31_7 <= 1'h0; // @[BitPlruReplacementPolicy.scala 87:45]
    end else if (5'h1f == io_control_setIdx) begin // @[BitPlruReplacementPolicy.scala 93:41]
      if (io_control_update_valid) begin // @[BitPlruReplacementPolicy.scala 96:37]
        REG_31_7 <= newMruBits_7; // @[BitPlruReplacementPolicy.scala 97:28]
      end
    end
    if (reset) begin // @[SharedCacheReplacementPolicyType.scala 40:30]
      replaceWayPipeReg <= 3'h0; // @[SharedCacheReplacementPolicyType.scala 40:30]
    end else if (_replaceWayPipeReg_T) begin // @[SharedCacheReplacementPolicyType.scala 41:14]
      if (_capacity_T_1[0]) begin // @[Mux.scala 47:70]
        replaceWayPipeReg <= 3'h0;
      end else if (_capacity_T_1[1]) begin // @[Mux.scala 47:70]
        replaceWayPipeReg <= 3'h1;
      end else begin
        replaceWayPipeReg <= _replaceWay_T_14;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG__0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG__1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG__2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG__3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG__4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG__5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG__6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG__7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_1_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_1_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_1_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG_1_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG_1_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  REG_1_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG_2_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG_2_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_2_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG_2_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG_2_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  REG_2_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  REG_2_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  REG_2_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG_3_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  REG_3_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  REG_3_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG_3_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  REG_3_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  REG_3_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  REG_3_6 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  REG_3_7 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  REG_4_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  REG_4_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  REG_4_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  REG_4_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  REG_4_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  REG_4_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  REG_4_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG_4_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG_5_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG_5_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG_5_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG_5_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG_5_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG_5_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_5_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG_5_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG_6_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG_6_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG_6_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG_6_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG_6_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  REG_6_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  REG_6_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  REG_6_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  REG_7_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  REG_7_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  REG_7_2 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  REG_7_3 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  REG_7_4 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  REG_7_5 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  REG_7_6 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  REG_7_7 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  REG_8_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  REG_8_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  REG_8_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  REG_8_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  REG_8_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  REG_8_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  REG_8_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  REG_8_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  REG_9_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  REG_9_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  REG_9_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  REG_9_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  REG_9_4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  REG_9_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  REG_9_6 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  REG_9_7 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  REG_10_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  REG_10_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  REG_10_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  REG_10_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  REG_10_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  REG_10_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  REG_10_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  REG_10_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  REG_11_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  REG_11_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG_11_2 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  REG_11_3 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  REG_11_4 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  REG_11_5 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  REG_11_6 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  REG_11_7 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  REG_12_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  REG_12_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  REG_12_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  REG_12_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG_12_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG_12_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  REG_12_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  REG_12_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG_13_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  REG_13_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  REG_13_2 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG_13_3 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG_13_4 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG_13_5 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  REG_13_6 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  REG_13_7 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG_14_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  REG_14_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG_14_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  REG_14_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  REG_14_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG_14_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG_14_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  REG_14_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG_15_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  REG_15_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  REG_15_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  REG_15_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  REG_15_4 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  REG_15_5 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  REG_15_6 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  REG_15_7 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  REG_16_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  REG_16_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  REG_16_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  REG_16_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  REG_16_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  REG_16_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  REG_16_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  REG_16_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  REG_17_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  REG_17_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  REG_17_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  REG_17_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  REG_17_4 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  REG_17_5 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  REG_17_6 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  REG_17_7 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  REG_18_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  REG_18_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  REG_18_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  REG_18_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  REG_18_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  REG_18_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  REG_18_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  REG_18_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  REG_19_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  REG_19_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  REG_19_2 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  REG_19_3 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  REG_19_4 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  REG_19_5 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  REG_19_6 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  REG_19_7 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  REG_20_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  REG_20_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  REG_20_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  REG_20_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  REG_20_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  REG_20_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  REG_20_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  REG_20_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  REG_21_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  REG_21_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  REG_21_2 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  REG_21_3 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  REG_21_4 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  REG_21_5 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  REG_21_6 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  REG_21_7 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  REG_22_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  REG_22_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  REG_22_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  REG_22_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  REG_22_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  REG_22_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  REG_22_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  REG_22_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  REG_23_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  REG_23_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  REG_23_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  REG_23_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  REG_23_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  REG_23_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  REG_23_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  REG_23_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  REG_24_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  REG_24_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  REG_24_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  REG_24_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  REG_24_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  REG_24_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  REG_24_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  REG_24_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  REG_25_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  REG_25_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  REG_25_2 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  REG_25_3 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  REG_25_4 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  REG_25_5 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  REG_25_6 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  REG_25_7 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  REG_26_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  REG_26_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  REG_26_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  REG_26_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  REG_26_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  REG_26_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  REG_26_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  REG_26_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  REG_27_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  REG_27_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  REG_27_2 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  REG_27_3 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  REG_27_4 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  REG_27_5 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  REG_27_6 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  REG_27_7 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  REG_28_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  REG_28_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  REG_28_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  REG_28_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  REG_28_4 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  REG_28_5 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  REG_28_6 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  REG_28_7 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  REG_29_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  REG_29_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  REG_29_2 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  REG_29_3 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  REG_29_4 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  REG_29_5 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  REG_29_6 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  REG_29_7 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  REG_30_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  REG_30_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  REG_30_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  REG_30_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  REG_30_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  REG_30_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  REG_30_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  REG_30_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  REG_31_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  REG_31_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  REG_31_2 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  REG_31_3 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  REG_31_4 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  REG_31_5 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  REG_31_6 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  REG_31_7 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  replaceWayPipeReg = _RAND_256[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SharedPipelinedCacheTop(
  input          clock,
  input          reset,
  output         io_cache_coreReqs_0_reqId_ready,
  input          io_cache_coreReqs_0_reqId_valid,
  input  [1:0]   io_cache_coreReqs_0_reqId_bits,
  input  [14:0]  io_cache_coreReqs_0_addr,
  input          io_cache_coreReqs_0_rw,
  input  [127:0] io_cache_coreReqs_0_wData,
  output         io_cache_coreReqs_1_reqId_ready,
  input          io_cache_coreReqs_1_reqId_valid,
  input  [1:0]   io_cache_coreReqs_1_reqId_bits,
  input  [14:0]  io_cache_coreReqs_1_addr,
  input          io_cache_coreReqs_1_rw,
  input  [127:0] io_cache_coreReqs_1_wData,
  output         io_cache_coreReqs_2_reqId_ready,
  input          io_cache_coreReqs_2_reqId_valid,
  input  [1:0]   io_cache_coreReqs_2_reqId_bits,
  input  [14:0]  io_cache_coreReqs_2_addr,
  input          io_cache_coreReqs_2_rw,
  input  [127:0] io_cache_coreReqs_2_wData,
  output         io_cache_coreReqs_3_reqId_ready,
  input          io_cache_coreReqs_3_reqId_valid,
  input  [1:0]   io_cache_coreReqs_3_reqId_bits,
  input  [14:0]  io_cache_coreReqs_3_addr,
  input          io_cache_coreReqs_3_rw,
  input  [127:0] io_cache_coreReqs_3_wData,
  output         io_cache_coreResps_0_reqId_valid,
  output [1:0]   io_cache_coreResps_0_reqId_bits,
  output [127:0] io_cache_coreResps_0_rData,
  output         io_cache_coreResps_0_responseStatus,
  output         io_cache_coreResps_1_reqId_valid,
  output [1:0]   io_cache_coreResps_1_reqId_bits,
  output [127:0] io_cache_coreResps_1_rData,
  output         io_cache_coreResps_1_responseStatus,
  output         io_cache_coreResps_2_reqId_valid,
  output [1:0]   io_cache_coreResps_2_reqId_bits,
  output [127:0] io_cache_coreResps_2_rData,
  output         io_cache_coreResps_2_responseStatus,
  output         io_cache_coreResps_3_reqId_valid,
  output [1:0]   io_cache_coreResps_3_reqId_bits,
  output [127:0] io_cache_coreResps_3_rData,
  output         io_cache_coreResps_3_responseStatus,
  input          io_mem_rChannel_rAddr_ready,
  output         io_mem_rChannel_rAddr_valid,
  output [14:0]  io_mem_rChannel_rAddr_bits,
  output         io_mem_rChannel_rData_ready,
  input          io_mem_rChannel_rData_valid,
  input  [15:0]  io_mem_rChannel_rData_bits,
  input          io_mem_rChannel_rLast,
  input          io_mem_wChannel_wAddr_ready,
  output         io_mem_wChannel_wAddr_valid,
  output [14:0]  io_mem_wChannel_wAddr_bits,
  input          io_mem_wChannel_wData_ready,
  output         io_mem_wChannel_wData_valid,
  output [15:0]  io_mem_wChannel_wData_bits,
  output         io_mem_wChannel_wLast
);
  wire  l2Cache_clock; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_reset; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_0_reqId_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_0_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreReqs_0_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [14:0] l2Cache_io_cache_coreReqs_0_addr; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_0_rw; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreReqs_0_wData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_1_reqId_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_1_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreReqs_1_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [14:0] l2Cache_io_cache_coreReqs_1_addr; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_1_rw; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreReqs_1_wData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_2_reqId_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_2_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreReqs_2_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [14:0] l2Cache_io_cache_coreReqs_2_addr; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_2_rw; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreReqs_2_wData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_3_reqId_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_3_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreReqs_3_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [14:0] l2Cache_io_cache_coreReqs_3_addr; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreReqs_3_rw; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreReqs_3_wData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_0_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreResps_0_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreResps_0_rData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_0_responseStatus; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_1_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreResps_1_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreResps_1_rData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_1_responseStatus; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_2_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreResps_2_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreResps_2_rData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_2_responseStatus; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_3_reqId_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [1:0] l2Cache_io_cache_coreResps_3_reqId_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [127:0] l2Cache_io_cache_coreResps_3_rData; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_cache_coreResps_3_responseStatus; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_repPol_update_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [2:0] l2Cache_io_repPol_update_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_repPol_stall; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [4:0] l2Cache_io_repPol_setIdx; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [2:0] l2Cache_io_repPol_replaceWay; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_rChannel_rAddr_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_rChannel_rAddr_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [14:0] l2Cache_io_mem_rChannel_rAddr_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_rChannel_rData_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_rChannel_rData_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [15:0] l2Cache_io_mem_rChannel_rData_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_rChannel_rLast; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_wChannel_wAddr_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_wChannel_wAddr_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [14:0] l2Cache_io_mem_wChannel_wAddr_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_wChannel_wData_ready; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_wChannel_wData_valid; // @[SharedPipelinedCacheTop.scala 28:23]
  wire [15:0] l2Cache_io_mem_wChannel_wData_bits; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  l2Cache_io_mem_wChannel_wLast; // @[SharedPipelinedCacheTop.scala 28:23]
  wire  repPol_clock; // @[SharedPipelinedCacheTop.scala 39:22]
  wire  repPol_reset; // @[SharedPipelinedCacheTop.scala 39:22]
  wire  repPol_io_control_update_valid; // @[SharedPipelinedCacheTop.scala 39:22]
  wire [2:0] repPol_io_control_update_bits; // @[SharedPipelinedCacheTop.scala 39:22]
  wire  repPol_io_control_stall; // @[SharedPipelinedCacheTop.scala 39:22]
  wire [4:0] repPol_io_control_setIdx; // @[SharedPipelinedCacheTop.scala 39:22]
  wire [2:0] repPol_io_control_replaceWay; // @[SharedPipelinedCacheTop.scala 39:22]
  SharedPipelinedCache l2Cache ( // @[SharedPipelinedCacheTop.scala 28:23]
    .clock(l2Cache_clock),
    .reset(l2Cache_reset),
    .io_cache_coreReqs_0_reqId_ready(l2Cache_io_cache_coreReqs_0_reqId_ready),
    .io_cache_coreReqs_0_reqId_valid(l2Cache_io_cache_coreReqs_0_reqId_valid),
    .io_cache_coreReqs_0_reqId_bits(l2Cache_io_cache_coreReqs_0_reqId_bits),
    .io_cache_coreReqs_0_addr(l2Cache_io_cache_coreReqs_0_addr),
    .io_cache_coreReqs_0_rw(l2Cache_io_cache_coreReqs_0_rw),
    .io_cache_coreReqs_0_wData(l2Cache_io_cache_coreReqs_0_wData),
    .io_cache_coreReqs_1_reqId_ready(l2Cache_io_cache_coreReqs_1_reqId_ready),
    .io_cache_coreReqs_1_reqId_valid(l2Cache_io_cache_coreReqs_1_reqId_valid),
    .io_cache_coreReqs_1_reqId_bits(l2Cache_io_cache_coreReqs_1_reqId_bits),
    .io_cache_coreReqs_1_addr(l2Cache_io_cache_coreReqs_1_addr),
    .io_cache_coreReqs_1_rw(l2Cache_io_cache_coreReqs_1_rw),
    .io_cache_coreReqs_1_wData(l2Cache_io_cache_coreReqs_1_wData),
    .io_cache_coreReqs_2_reqId_ready(l2Cache_io_cache_coreReqs_2_reqId_ready),
    .io_cache_coreReqs_2_reqId_valid(l2Cache_io_cache_coreReqs_2_reqId_valid),
    .io_cache_coreReqs_2_reqId_bits(l2Cache_io_cache_coreReqs_2_reqId_bits),
    .io_cache_coreReqs_2_addr(l2Cache_io_cache_coreReqs_2_addr),
    .io_cache_coreReqs_2_rw(l2Cache_io_cache_coreReqs_2_rw),
    .io_cache_coreReqs_2_wData(l2Cache_io_cache_coreReqs_2_wData),
    .io_cache_coreReqs_3_reqId_ready(l2Cache_io_cache_coreReqs_3_reqId_ready),
    .io_cache_coreReqs_3_reqId_valid(l2Cache_io_cache_coreReqs_3_reqId_valid),
    .io_cache_coreReqs_3_reqId_bits(l2Cache_io_cache_coreReqs_3_reqId_bits),
    .io_cache_coreReqs_3_addr(l2Cache_io_cache_coreReqs_3_addr),
    .io_cache_coreReqs_3_rw(l2Cache_io_cache_coreReqs_3_rw),
    .io_cache_coreReqs_3_wData(l2Cache_io_cache_coreReqs_3_wData),
    .io_cache_coreResps_0_reqId_valid(l2Cache_io_cache_coreResps_0_reqId_valid),
    .io_cache_coreResps_0_reqId_bits(l2Cache_io_cache_coreResps_0_reqId_bits),
    .io_cache_coreResps_0_rData(l2Cache_io_cache_coreResps_0_rData),
    .io_cache_coreResps_0_responseStatus(l2Cache_io_cache_coreResps_0_responseStatus),
    .io_cache_coreResps_1_reqId_valid(l2Cache_io_cache_coreResps_1_reqId_valid),
    .io_cache_coreResps_1_reqId_bits(l2Cache_io_cache_coreResps_1_reqId_bits),
    .io_cache_coreResps_1_rData(l2Cache_io_cache_coreResps_1_rData),
    .io_cache_coreResps_1_responseStatus(l2Cache_io_cache_coreResps_1_responseStatus),
    .io_cache_coreResps_2_reqId_valid(l2Cache_io_cache_coreResps_2_reqId_valid),
    .io_cache_coreResps_2_reqId_bits(l2Cache_io_cache_coreResps_2_reqId_bits),
    .io_cache_coreResps_2_rData(l2Cache_io_cache_coreResps_2_rData),
    .io_cache_coreResps_2_responseStatus(l2Cache_io_cache_coreResps_2_responseStatus),
    .io_cache_coreResps_3_reqId_valid(l2Cache_io_cache_coreResps_3_reqId_valid),
    .io_cache_coreResps_3_reqId_bits(l2Cache_io_cache_coreResps_3_reqId_bits),
    .io_cache_coreResps_3_rData(l2Cache_io_cache_coreResps_3_rData),
    .io_cache_coreResps_3_responseStatus(l2Cache_io_cache_coreResps_3_responseStatus),
    .io_repPol_update_valid(l2Cache_io_repPol_update_valid),
    .io_repPol_update_bits(l2Cache_io_repPol_update_bits),
    .io_repPol_stall(l2Cache_io_repPol_stall),
    .io_repPol_setIdx(l2Cache_io_repPol_setIdx),
    .io_repPol_replaceWay(l2Cache_io_repPol_replaceWay),
    .io_mem_rChannel_rAddr_ready(l2Cache_io_mem_rChannel_rAddr_ready),
    .io_mem_rChannel_rAddr_valid(l2Cache_io_mem_rChannel_rAddr_valid),
    .io_mem_rChannel_rAddr_bits(l2Cache_io_mem_rChannel_rAddr_bits),
    .io_mem_rChannel_rData_ready(l2Cache_io_mem_rChannel_rData_ready),
    .io_mem_rChannel_rData_valid(l2Cache_io_mem_rChannel_rData_valid),
    .io_mem_rChannel_rData_bits(l2Cache_io_mem_rChannel_rData_bits),
    .io_mem_rChannel_rLast(l2Cache_io_mem_rChannel_rLast),
    .io_mem_wChannel_wAddr_ready(l2Cache_io_mem_wChannel_wAddr_ready),
    .io_mem_wChannel_wAddr_valid(l2Cache_io_mem_wChannel_wAddr_valid),
    .io_mem_wChannel_wAddr_bits(l2Cache_io_mem_wChannel_wAddr_bits),
    .io_mem_wChannel_wData_ready(l2Cache_io_mem_wChannel_wData_ready),
    .io_mem_wChannel_wData_valid(l2Cache_io_mem_wChannel_wData_valid),
    .io_mem_wChannel_wData_bits(l2Cache_io_mem_wChannel_wData_bits),
    .io_mem_wChannel_wLast(l2Cache_io_mem_wChannel_wLast)
  );
  BitPlruReplacementPolicy repPol ( // @[SharedPipelinedCacheTop.scala 39:22]
    .clock(repPol_clock),
    .reset(repPol_reset),
    .io_control_update_valid(repPol_io_control_update_valid),
    .io_control_update_bits(repPol_io_control_update_bits),
    .io_control_stall(repPol_io_control_stall),
    .io_control_setIdx(repPol_io_control_setIdx),
    .io_control_replaceWay(repPol_io_control_replaceWay)
  );
  assign io_cache_coreReqs_0_reqId_ready = l2Cache_io_cache_coreReqs_0_reqId_ready; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreReqs_1_reqId_ready = l2Cache_io_cache_coreReqs_1_reqId_ready; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreReqs_2_reqId_ready = l2Cache_io_cache_coreReqs_2_reqId_ready; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreReqs_3_reqId_ready = l2Cache_io_cache_coreReqs_3_reqId_ready; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_0_reqId_valid = l2Cache_io_cache_coreResps_0_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_0_reqId_bits = l2Cache_io_cache_coreResps_0_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_0_rData = l2Cache_io_cache_coreResps_0_rData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_0_responseStatus = l2Cache_io_cache_coreResps_0_responseStatus; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_1_reqId_valid = l2Cache_io_cache_coreResps_1_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_1_reqId_bits = l2Cache_io_cache_coreResps_1_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_1_rData = l2Cache_io_cache_coreResps_1_rData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_1_responseStatus = l2Cache_io_cache_coreResps_1_responseStatus; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_2_reqId_valid = l2Cache_io_cache_coreResps_2_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_2_reqId_bits = l2Cache_io_cache_coreResps_2_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_2_rData = l2Cache_io_cache_coreResps_2_rData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_2_responseStatus = l2Cache_io_cache_coreResps_2_responseStatus; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_3_reqId_valid = l2Cache_io_cache_coreResps_3_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_3_reqId_bits = l2Cache_io_cache_coreResps_3_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_3_rData = l2Cache_io_cache_coreResps_3_rData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_cache_coreResps_3_responseStatus = l2Cache_io_cache_coreResps_3_responseStatus; // @[SharedPipelinedCacheTop.scala 43:20]
  assign io_mem_rChannel_rAddr_valid = l2Cache_io_mem_rChannel_rAddr_valid; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_rChannel_rAddr_bits = l2Cache_io_mem_rChannel_rAddr_bits; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_rChannel_rData_ready = l2Cache_io_mem_rChannel_rData_ready; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_wChannel_wAddr_valid = l2Cache_io_mem_wChannel_wAddr_valid; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_wChannel_wAddr_bits = l2Cache_io_mem_wChannel_wAddr_bits; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_wChannel_wData_valid = l2Cache_io_mem_wChannel_wData_valid; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_wChannel_wData_bits = l2Cache_io_mem_wChannel_wData_bits; // @[SharedPipelinedCacheTop.scala 44:18]
  assign io_mem_wChannel_wLast = l2Cache_io_mem_wChannel_wLast; // @[SharedPipelinedCacheTop.scala 44:18]
  assign l2Cache_clock = clock;
  assign l2Cache_reset = reset;
  assign l2Cache_io_cache_coreReqs_0_reqId_valid = io_cache_coreReqs_0_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_0_reqId_bits = io_cache_coreReqs_0_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_0_addr = io_cache_coreReqs_0_addr; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_0_rw = io_cache_coreReqs_0_rw; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_0_wData = io_cache_coreReqs_0_wData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_1_reqId_valid = io_cache_coreReqs_1_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_1_reqId_bits = io_cache_coreReqs_1_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_1_addr = io_cache_coreReqs_1_addr; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_1_rw = io_cache_coreReqs_1_rw; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_1_wData = io_cache_coreReqs_1_wData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_2_reqId_valid = io_cache_coreReqs_2_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_2_reqId_bits = io_cache_coreReqs_2_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_2_addr = io_cache_coreReqs_2_addr; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_2_rw = io_cache_coreReqs_2_rw; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_2_wData = io_cache_coreReqs_2_wData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_3_reqId_valid = io_cache_coreReqs_3_reqId_valid; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_3_reqId_bits = io_cache_coreReqs_3_reqId_bits; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_3_addr = io_cache_coreReqs_3_addr; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_3_rw = io_cache_coreReqs_3_rw; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_cache_coreReqs_3_wData = io_cache_coreReqs_3_wData; // @[SharedPipelinedCacheTop.scala 43:20]
  assign l2Cache_io_repPol_replaceWay = repPol_io_control_replaceWay; // @[SharedPipelinedCacheTop.scala 42:21]
  assign l2Cache_io_mem_rChannel_rAddr_ready = io_mem_rChannel_rAddr_ready; // @[SharedPipelinedCacheTop.scala 44:18]
  assign l2Cache_io_mem_rChannel_rData_valid = io_mem_rChannel_rData_valid; // @[SharedPipelinedCacheTop.scala 44:18]
  assign l2Cache_io_mem_rChannel_rData_bits = io_mem_rChannel_rData_bits; // @[SharedPipelinedCacheTop.scala 44:18]
  assign l2Cache_io_mem_rChannel_rLast = io_mem_rChannel_rLast; // @[SharedPipelinedCacheTop.scala 44:18]
  assign l2Cache_io_mem_wChannel_wAddr_ready = io_mem_wChannel_wAddr_ready; // @[SharedPipelinedCacheTop.scala 44:18]
  assign l2Cache_io_mem_wChannel_wData_ready = io_mem_wChannel_wData_ready; // @[SharedPipelinedCacheTop.scala 44:18]
  assign repPol_clock = clock;
  assign repPol_reset = reset;
  assign repPol_io_control_update_valid = l2Cache_io_repPol_update_valid; // @[SharedPipelinedCacheTop.scala 42:21]
  assign repPol_io_control_update_bits = l2Cache_io_repPol_update_bits; // @[SharedPipelinedCacheTop.scala 42:21]
  assign repPol_io_control_stall = l2Cache_io_repPol_stall; // @[SharedPipelinedCacheTop.scala 42:21]
  assign repPol_io_control_setIdx = l2Cache_io_repPol_setIdx; // @[SharedPipelinedCacheTop.scala 42:21]
endmodule
module MemBlock_40(
  input         clock,
  input  [13:0] io_readAddr,
  input  [13:0] io_writeAddr,
  input  [15:0] io_writeData,
  input         io_wrEn,
  output [15:0] io_readData
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] mem [0:16383]; // @[MemBlock.scala 29:24]
  wire  mem_readData_MPORT_en; // @[MemBlock.scala 29:24]
  wire [13:0] mem_readData_MPORT_addr; // @[MemBlock.scala 29:24]
  wire [15:0] mem_readData_MPORT_data; // @[MemBlock.scala 29:24]
  wire [15:0] mem_MPORT_data; // @[MemBlock.scala 29:24]
  wire [13:0] mem_MPORT_addr; // @[MemBlock.scala 29:24]
  wire  mem_MPORT_mask; // @[MemBlock.scala 29:24]
  wire  mem_MPORT_en; // @[MemBlock.scala 29:24]
  reg [15:0] mem_readData_MPORT_data_pipe_0;
  reg [15:0] writeDataReg; // @[MemBlock.scala 50:29]
  reg  forwardSelReg; // @[MemBlock.scala 51:30]
  wire [15:0] readData = mem_readData_MPORT_data_pipe_0; // @[MemBlock.scala 28:29 48:12]
  assign mem_readData_MPORT_en = 1'h1;
  assign mem_readData_MPORT_addr = io_readAddr;
  assign mem_readData_MPORT_data = mem[mem_readData_MPORT_addr]; // @[MemBlock.scala 29:24]
  assign mem_MPORT_data = io_writeData;
  assign mem_MPORT_addr = io_writeAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEn;
  assign io_readData = forwardSelReg ? writeDataReg : readData; // @[MemBlock.scala 52:21]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[MemBlock.scala 29:24]
    end
    if (1'h1) begin
      mem_readData_MPORT_data_pipe_0 <= mem_readData_MPORT_data;
    end
    writeDataReg <= io_writeData; // @[MemBlock.scala 50:29]
    forwardSelReg <= io_writeAddr == io_readAddr & io_wrEn; // @[MemBlock.scala 51:62]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
  integer initvar;
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_readData_MPORT_data_pipe_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  writeDataReg = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  forwardSelReg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
  $readmemh("test_mem_32w.hex", mem);
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyMemory(
  input         clock,
  input         reset,
  output        io_rChannel_rAddr_ready,
  input         io_rChannel_rAddr_valid,
  input  [13:0] io_rChannel_rAddr_bits,
  input         io_rChannel_rData_ready,
  output        io_rChannel_rData_valid,
  output [15:0] io_rChannel_rData_bits,
  output        io_rChannel_rLast,
  output        io_wChannel_wAddr_ready,
  input         io_wChannel_wAddr_valid,
  input  [13:0] io_wChannel_wAddr_bits,
  output        io_wChannel_wData_ready,
  input         io_wChannel_wData_valid,
  input  [15:0] io_wChannel_wData_bits,
  input         io_wChannel_wLast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  mem_clock; // @[DummyMemory.scala 32:19]
  wire [13:0] mem_io_readAddr; // @[DummyMemory.scala 32:19]
  wire [13:0] mem_io_writeAddr; // @[DummyMemory.scala 32:19]
  wire [15:0] mem_io_writeData; // @[DummyMemory.scala 32:19]
  wire  mem_io_wrEn; // @[DummyMemory.scala 32:19]
  wire [15:0] mem_io_readData; // @[DummyMemory.scala 32:19]
  reg [1:0] stateReg; // @[DummyMemory.scala 16:25]
  reg [13:0] addrReg; // @[DummyMemory.scala 17:24]
  reg [4:0] burstCountReg; // @[DummyMemory.scala 18:30]
  wire  rAddrReady = 2'h0 == stateReg; // @[DummyMemory.scala 39:20]
  wire [13:0] _GEN_2 = io_rChannel_rAddr_valid ? io_rChannel_rAddr_bits : 14'h0; // @[DummyMemory.scala 44:37 45:21 27:32]
  wire [4:0] _nextBurstCount_T_1 = burstCountReg + 5'h1; // @[DummyMemory.scala 62:41]
  wire [13:0] _nextReadAddr_T_1 = addrReg + 14'h1; // @[DummyMemory.scala 63:33]
  wire  _T_2 = burstCountReg == 5'h1f; // @[DummyMemory.scala 65:28]
  wire [1:0] _GEN_6 = burstCountReg == 5'h1f ? 2'h0 : stateReg; // @[DummyMemory.scala 65:49 67:20 16:25]
  wire [4:0] _GEN_7 = burstCountReg == 5'h1f ? 5'h0 : _nextBurstCount_T_1; // @[DummyMemory.scala 62:24 65:49 68:26]
  wire [13:0] nextReadAddr = burstCountReg == 5'h1f ? 14'h0 : _nextReadAddr_T_1; // @[DummyMemory.scala 63:22 65:49 69:24]
  wire  _GEN_9 = io_rChannel_rData_ready & _T_2; // @[DummyMemory.scala 24:26 59:37]
  wire [13:0] _GEN_11 = io_rChannel_rData_ready ? nextReadAddr : addrReg; // @[DummyMemory.scala 57:19 59:37 72:21]
  wire [31:0] nextBurstCount = {{27'd0}, _GEN_7}; // @[DummyMemory.scala 61:41]
  wire [31:0] _GEN_12 = io_rChannel_rData_ready ? nextBurstCount : {{27'd0}, burstCountReg}; // @[DummyMemory.scala 59:37 74:23 18:30]
  wire [1:0] _GEN_13 = io_wChannel_wLast | _T_2 ? 2'h0 : stateReg; // @[DummyMemory.scala 91:70 92:20 16:25]
  wire [4:0] _GEN_14 = io_wChannel_wLast | _T_2 ? 5'h0 : _nextBurstCount_T_1; // @[DummyMemory.scala 87:24 91:70 93:26]
  wire [13:0] nextWriteAddr = io_wChannel_wLast | _T_2 ? 14'h0 : _nextReadAddr_T_1; // @[DummyMemory.scala 86:23 91:70 94:25]
  wire [15:0] _GEN_16 = io_wChannel_wData_valid ? 16'h1 : 16'h0; // @[DummyMemory.scala 83:37 89:17 30:28]
  wire [1:0] _GEN_17 = io_wChannel_wData_valid ? _GEN_13 : stateReg; // @[DummyMemory.scala 16:25 83:37]
  wire [13:0] _GEN_18 = io_wChannel_wData_valid ? nextWriteAddr : addrReg; // @[DummyMemory.scala 83:37 97:17 17:24]
  wire [31:0] nextBurstCount_1 = {{27'd0}, _GEN_14}; // @[DummyMemory.scala 85:41]
  wire [31:0] _GEN_19 = io_wChannel_wData_valid ? nextBurstCount_1 : {{27'd0}, burstCountReg}; // @[DummyMemory.scala 83:37 98:23 18:30]
  wire [13:0] _GEN_21 = 2'h2 == stateReg ? addrReg : 14'h0; // @[DummyMemory.scala 39:20 80:20 28:33]
  wire [15:0] _GEN_22 = 2'h2 == stateReg ? io_wChannel_wData_bits : 16'h0; // @[DummyMemory.scala 39:20 81:20 29:33]
  wire [15:0] _GEN_23 = 2'h2 == stateReg ? _GEN_16 : 16'h0; // @[DummyMemory.scala 39:20 30:28]
  wire [31:0] _GEN_26 = 2'h2 == stateReg ? _GEN_19 : {{27'd0}, burstCountReg}; // @[DummyMemory.scala 39:20 18:30]
  wire [15:0] _GEN_27 = 2'h1 == stateReg ? mem_io_readData : 16'h0; // @[DummyMemory.scala 39:20 55:17 23:30]
  wire [13:0] _GEN_29 = 2'h1 == stateReg ? _GEN_11 : 14'h0; // @[DummyMemory.scala 39:20 27:32]
  wire [31:0] _GEN_33 = 2'h1 == stateReg ? _GEN_12 : _GEN_26; // @[DummyMemory.scala 39:20]
  wire  _GEN_34 = 2'h1 == stateReg ? 1'h0 : 2'h2 == stateReg; // @[DummyMemory.scala 39:20 26:31]
  wire [13:0] _GEN_35 = 2'h1 == stateReg ? 14'h0 : _GEN_21; // @[DummyMemory.scala 39:20 28:33]
  wire [15:0] _GEN_36 = 2'h1 == stateReg ? 16'h0 : _GEN_22; // @[DummyMemory.scala 39:20 29:33]
  wire [15:0] _GEN_37 = 2'h1 == stateReg ? 16'h0 : _GEN_23; // @[DummyMemory.scala 39:20 30:28]
  wire [31:0] _GEN_45 = rAddrReady ? {{27'd0}, burstCountReg} : _GEN_33; // @[DummyMemory.scala 39:20 18:30]
  wire [15:0] memWrEn = rAddrReady ? 16'h0 : _GEN_37; // @[DummyMemory.scala 39:20 30:28]
  wire [31:0] _GEN_50 = reset ? 32'h0 : _GEN_45; // @[DummyMemory.scala 18:{30,30}]
  MemBlock_40 mem ( // @[DummyMemory.scala 32:19]
    .clock(mem_clock),
    .io_readAddr(mem_io_readAddr),
    .io_writeAddr(mem_io_writeAddr),
    .io_writeData(mem_io_writeData),
    .io_wrEn(mem_io_wrEn),
    .io_readData(mem_io_readData)
  );
  assign io_rChannel_rAddr_ready = 2'h0 == stateReg; // @[DummyMemory.scala 39:20]
  assign io_rChannel_rData_valid = rAddrReady ? 1'h0 : 2'h1 == stateReg; // @[DummyMemory.scala 39:20 22:31]
  assign io_rChannel_rData_bits = rAddrReady ? 16'h0 : _GEN_27; // @[DummyMemory.scala 39:20 23:30]
  assign io_rChannel_rLast = rAddrReady ? 1'h0 : 2'h1 == stateReg & _GEN_9; // @[DummyMemory.scala 39:20 24:26]
  assign io_wChannel_wAddr_ready = 2'h0 == stateReg; // @[DummyMemory.scala 39:20]
  assign io_wChannel_wData_ready = rAddrReady ? 1'h0 : _GEN_34; // @[DummyMemory.scala 39:20 26:31]
  assign mem_clock = clock;
  assign mem_io_readAddr = rAddrReady ? _GEN_2 : _GEN_29; // @[DummyMemory.scala 39:20]
  assign mem_io_writeAddr = rAddrReady ? 14'h0 : _GEN_35; // @[DummyMemory.scala 39:20 28:33]
  assign mem_io_writeData = rAddrReady ? 16'h0 : _GEN_36; // @[DummyMemory.scala 39:20 29:33]
  assign mem_io_wrEn = memWrEn[0]; // @[DummyMemory.scala 37:15]
  always @(posedge clock) begin
    if (reset) begin // @[DummyMemory.scala 16:25]
      stateReg <= 2'h0; // @[DummyMemory.scala 16:25]
    end else if (rAddrReady) begin // @[DummyMemory.scala 39:20]
      if (io_rChannel_rAddr_valid) begin // @[DummyMemory.scala 44:37]
        stateReg <= 2'h1; // @[DummyMemory.scala 47:18]
      end else if (io_wChannel_wAddr_valid) begin // @[DummyMemory.scala 48:44]
        stateReg <= 2'h2; // @[DummyMemory.scala 50:18]
      end
    end else if (2'h1 == stateReg) begin // @[DummyMemory.scala 39:20]
      if (io_rChannel_rData_ready) begin // @[DummyMemory.scala 59:37]
        stateReg <= _GEN_6;
      end
    end else if (2'h2 == stateReg) begin // @[DummyMemory.scala 39:20]
      stateReg <= _GEN_17;
    end
    if (reset) begin // @[DummyMemory.scala 17:24]
      addrReg <= 14'h0; // @[DummyMemory.scala 17:24]
    end else if (rAddrReady) begin // @[DummyMemory.scala 39:20]
      if (io_rChannel_rAddr_valid) begin // @[DummyMemory.scala 44:37]
        addrReg <= io_rChannel_rAddr_bits; // @[DummyMemory.scala 46:17]
      end else if (io_wChannel_wAddr_valid) begin // @[DummyMemory.scala 48:44]
        addrReg <= io_wChannel_wAddr_bits; // @[DummyMemory.scala 49:17]
      end
    end else if (2'h1 == stateReg) begin // @[DummyMemory.scala 39:20]
      if (io_rChannel_rData_ready) begin // @[DummyMemory.scala 59:37]
        addrReg <= nextReadAddr; // @[DummyMemory.scala 72:21]
      end
    end else if (2'h2 == stateReg) begin // @[DummyMemory.scala 39:20]
      addrReg <= _GEN_18;
    end
    burstCountReg <= _GEN_50[4:0]; // @[DummyMemory.scala 18:{30,30}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  addrReg = _RAND_1[13:0];
  _RAND_2 = {1{`RANDOM}};
  burstCountReg = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SharedPipelinedCacheTestTopDe2115(
  input         clock,
  input         reset,
  input         io_rxd,
  output        io_txd,
  input         io_scheduler_coreId_valid,
  input  [1:0]  io_scheduler_coreId_bits,
  input         io_scheduler_setCritical,
  input         io_scheduler_unsetCritical,
  input  [10:0] io_scheduler_contentionLimit
);
  wire  cacheReqCtrl_clock; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_reset; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_rxd; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_txd; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_0_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_0_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreReqs_0_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [14:0] cacheReqCtrl_io_cache_coreReqs_0_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_0_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreReqs_0_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_1_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_1_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreReqs_1_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [14:0] cacheReqCtrl_io_cache_coreReqs_1_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_1_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreReqs_1_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_2_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_2_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreReqs_2_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [14:0] cacheReqCtrl_io_cache_coreReqs_2_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_2_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreReqs_2_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_3_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_3_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreReqs_3_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [14:0] cacheReqCtrl_io_cache_coreReqs_3_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreReqs_3_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreReqs_3_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_0_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreResps_0_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreResps_0_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_0_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_1_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreResps_1_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreResps_1_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_1_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_2_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreResps_2_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreResps_2_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_2_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_3_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [1:0] cacheReqCtrl_io_cache_coreResps_3_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire [127:0] cacheReqCtrl_io_cache_coreResps_3_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  cacheReqCtrl_io_cache_coreResps_3_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
  wire  l2Cache_clock; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_reset; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_0_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_0_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreReqs_0_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [14:0] l2Cache_io_cache_coreReqs_0_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_0_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreReqs_0_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_1_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_1_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreReqs_1_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [14:0] l2Cache_io_cache_coreReqs_1_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_1_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreReqs_1_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_2_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_2_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreReqs_2_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [14:0] l2Cache_io_cache_coreReqs_2_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_2_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreReqs_2_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_3_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_3_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreReqs_3_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [14:0] l2Cache_io_cache_coreReqs_3_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreReqs_3_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreReqs_3_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_0_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreResps_0_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreResps_0_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_0_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_1_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreResps_1_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreResps_1_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_1_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_2_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreResps_2_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreResps_2_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_2_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_3_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [1:0] l2Cache_io_cache_coreResps_3_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [127:0] l2Cache_io_cache_coreResps_3_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_cache_coreResps_3_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_rChannel_rAddr_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_rChannel_rAddr_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [14:0] l2Cache_io_mem_rChannel_rAddr_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_rChannel_rData_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_rChannel_rData_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [15:0] l2Cache_io_mem_rChannel_rData_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_rChannel_rLast; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_wChannel_wAddr_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_wChannel_wAddr_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [14:0] l2Cache_io_mem_wChannel_wAddr_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_wChannel_wData_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_wChannel_wData_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire [15:0] l2Cache_io_mem_wChannel_wData_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  l2Cache_io_mem_wChannel_wLast; // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
  wire  memory_clock; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_reset; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_rChannel_rAddr_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_rChannel_rAddr_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire [13:0] memory_io_rChannel_rAddr_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_rChannel_rData_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_rChannel_rData_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire [15:0] memory_io_rChannel_rData_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_rChannel_rLast; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_wChannel_wAddr_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_wChannel_wAddr_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire [13:0] memory_io_wChannel_wAddr_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_wChannel_wData_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_wChannel_wData_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire [15:0] memory_io_wChannel_wData_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  wire  memory_io_wChannel_wLast; // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
  CacheRequestController cacheReqCtrl ( // @[SharedPipelinedCacheTestTopDe2115.scala 36:28]
    .clock(cacheReqCtrl_clock),
    .reset(cacheReqCtrl_reset),
    .io_rxd(cacheReqCtrl_io_rxd),
    .io_txd(cacheReqCtrl_io_txd),
    .io_cache_coreReqs_0_reqId_ready(cacheReqCtrl_io_cache_coreReqs_0_reqId_ready),
    .io_cache_coreReqs_0_reqId_valid(cacheReqCtrl_io_cache_coreReqs_0_reqId_valid),
    .io_cache_coreReqs_0_reqId_bits(cacheReqCtrl_io_cache_coreReqs_0_reqId_bits),
    .io_cache_coreReqs_0_addr(cacheReqCtrl_io_cache_coreReqs_0_addr),
    .io_cache_coreReqs_0_rw(cacheReqCtrl_io_cache_coreReqs_0_rw),
    .io_cache_coreReqs_0_wData(cacheReqCtrl_io_cache_coreReqs_0_wData),
    .io_cache_coreReqs_1_reqId_ready(cacheReqCtrl_io_cache_coreReqs_1_reqId_ready),
    .io_cache_coreReqs_1_reqId_valid(cacheReqCtrl_io_cache_coreReqs_1_reqId_valid),
    .io_cache_coreReqs_1_reqId_bits(cacheReqCtrl_io_cache_coreReqs_1_reqId_bits),
    .io_cache_coreReqs_1_addr(cacheReqCtrl_io_cache_coreReqs_1_addr),
    .io_cache_coreReqs_1_rw(cacheReqCtrl_io_cache_coreReqs_1_rw),
    .io_cache_coreReqs_1_wData(cacheReqCtrl_io_cache_coreReqs_1_wData),
    .io_cache_coreReqs_2_reqId_ready(cacheReqCtrl_io_cache_coreReqs_2_reqId_ready),
    .io_cache_coreReqs_2_reqId_valid(cacheReqCtrl_io_cache_coreReqs_2_reqId_valid),
    .io_cache_coreReqs_2_reqId_bits(cacheReqCtrl_io_cache_coreReqs_2_reqId_bits),
    .io_cache_coreReqs_2_addr(cacheReqCtrl_io_cache_coreReqs_2_addr),
    .io_cache_coreReqs_2_rw(cacheReqCtrl_io_cache_coreReqs_2_rw),
    .io_cache_coreReqs_2_wData(cacheReqCtrl_io_cache_coreReqs_2_wData),
    .io_cache_coreReqs_3_reqId_ready(cacheReqCtrl_io_cache_coreReqs_3_reqId_ready),
    .io_cache_coreReqs_3_reqId_valid(cacheReqCtrl_io_cache_coreReqs_3_reqId_valid),
    .io_cache_coreReqs_3_reqId_bits(cacheReqCtrl_io_cache_coreReqs_3_reqId_bits),
    .io_cache_coreReqs_3_addr(cacheReqCtrl_io_cache_coreReqs_3_addr),
    .io_cache_coreReqs_3_rw(cacheReqCtrl_io_cache_coreReqs_3_rw),
    .io_cache_coreReqs_3_wData(cacheReqCtrl_io_cache_coreReqs_3_wData),
    .io_cache_coreResps_0_reqId_valid(cacheReqCtrl_io_cache_coreResps_0_reqId_valid),
    .io_cache_coreResps_0_reqId_bits(cacheReqCtrl_io_cache_coreResps_0_reqId_bits),
    .io_cache_coreResps_0_rData(cacheReqCtrl_io_cache_coreResps_0_rData),
    .io_cache_coreResps_0_responseStatus(cacheReqCtrl_io_cache_coreResps_0_responseStatus),
    .io_cache_coreResps_1_reqId_valid(cacheReqCtrl_io_cache_coreResps_1_reqId_valid),
    .io_cache_coreResps_1_reqId_bits(cacheReqCtrl_io_cache_coreResps_1_reqId_bits),
    .io_cache_coreResps_1_rData(cacheReqCtrl_io_cache_coreResps_1_rData),
    .io_cache_coreResps_1_responseStatus(cacheReqCtrl_io_cache_coreResps_1_responseStatus),
    .io_cache_coreResps_2_reqId_valid(cacheReqCtrl_io_cache_coreResps_2_reqId_valid),
    .io_cache_coreResps_2_reqId_bits(cacheReqCtrl_io_cache_coreResps_2_reqId_bits),
    .io_cache_coreResps_2_rData(cacheReqCtrl_io_cache_coreResps_2_rData),
    .io_cache_coreResps_2_responseStatus(cacheReqCtrl_io_cache_coreResps_2_responseStatus),
    .io_cache_coreResps_3_reqId_valid(cacheReqCtrl_io_cache_coreResps_3_reqId_valid),
    .io_cache_coreResps_3_reqId_bits(cacheReqCtrl_io_cache_coreResps_3_reqId_bits),
    .io_cache_coreResps_3_rData(cacheReqCtrl_io_cache_coreResps_3_rData),
    .io_cache_coreResps_3_responseStatus(cacheReqCtrl_io_cache_coreResps_3_responseStatus)
  );
  SharedPipelinedCacheTop l2Cache ( // @[SharedPipelinedCacheTestTopDe2115.scala 38:23]
    .clock(l2Cache_clock),
    .reset(l2Cache_reset),
    .io_cache_coreReqs_0_reqId_ready(l2Cache_io_cache_coreReqs_0_reqId_ready),
    .io_cache_coreReqs_0_reqId_valid(l2Cache_io_cache_coreReqs_0_reqId_valid),
    .io_cache_coreReqs_0_reqId_bits(l2Cache_io_cache_coreReqs_0_reqId_bits),
    .io_cache_coreReqs_0_addr(l2Cache_io_cache_coreReqs_0_addr),
    .io_cache_coreReqs_0_rw(l2Cache_io_cache_coreReqs_0_rw),
    .io_cache_coreReqs_0_wData(l2Cache_io_cache_coreReqs_0_wData),
    .io_cache_coreReqs_1_reqId_ready(l2Cache_io_cache_coreReqs_1_reqId_ready),
    .io_cache_coreReqs_1_reqId_valid(l2Cache_io_cache_coreReqs_1_reqId_valid),
    .io_cache_coreReqs_1_reqId_bits(l2Cache_io_cache_coreReqs_1_reqId_bits),
    .io_cache_coreReqs_1_addr(l2Cache_io_cache_coreReqs_1_addr),
    .io_cache_coreReqs_1_rw(l2Cache_io_cache_coreReqs_1_rw),
    .io_cache_coreReqs_1_wData(l2Cache_io_cache_coreReqs_1_wData),
    .io_cache_coreReqs_2_reqId_ready(l2Cache_io_cache_coreReqs_2_reqId_ready),
    .io_cache_coreReqs_2_reqId_valid(l2Cache_io_cache_coreReqs_2_reqId_valid),
    .io_cache_coreReqs_2_reqId_bits(l2Cache_io_cache_coreReqs_2_reqId_bits),
    .io_cache_coreReqs_2_addr(l2Cache_io_cache_coreReqs_2_addr),
    .io_cache_coreReqs_2_rw(l2Cache_io_cache_coreReqs_2_rw),
    .io_cache_coreReqs_2_wData(l2Cache_io_cache_coreReqs_2_wData),
    .io_cache_coreReqs_3_reqId_ready(l2Cache_io_cache_coreReqs_3_reqId_ready),
    .io_cache_coreReqs_3_reqId_valid(l2Cache_io_cache_coreReqs_3_reqId_valid),
    .io_cache_coreReqs_3_reqId_bits(l2Cache_io_cache_coreReqs_3_reqId_bits),
    .io_cache_coreReqs_3_addr(l2Cache_io_cache_coreReqs_3_addr),
    .io_cache_coreReqs_3_rw(l2Cache_io_cache_coreReqs_3_rw),
    .io_cache_coreReqs_3_wData(l2Cache_io_cache_coreReqs_3_wData),
    .io_cache_coreResps_0_reqId_valid(l2Cache_io_cache_coreResps_0_reqId_valid),
    .io_cache_coreResps_0_reqId_bits(l2Cache_io_cache_coreResps_0_reqId_bits),
    .io_cache_coreResps_0_rData(l2Cache_io_cache_coreResps_0_rData),
    .io_cache_coreResps_0_responseStatus(l2Cache_io_cache_coreResps_0_responseStatus),
    .io_cache_coreResps_1_reqId_valid(l2Cache_io_cache_coreResps_1_reqId_valid),
    .io_cache_coreResps_1_reqId_bits(l2Cache_io_cache_coreResps_1_reqId_bits),
    .io_cache_coreResps_1_rData(l2Cache_io_cache_coreResps_1_rData),
    .io_cache_coreResps_1_responseStatus(l2Cache_io_cache_coreResps_1_responseStatus),
    .io_cache_coreResps_2_reqId_valid(l2Cache_io_cache_coreResps_2_reqId_valid),
    .io_cache_coreResps_2_reqId_bits(l2Cache_io_cache_coreResps_2_reqId_bits),
    .io_cache_coreResps_2_rData(l2Cache_io_cache_coreResps_2_rData),
    .io_cache_coreResps_2_responseStatus(l2Cache_io_cache_coreResps_2_responseStatus),
    .io_cache_coreResps_3_reqId_valid(l2Cache_io_cache_coreResps_3_reqId_valid),
    .io_cache_coreResps_3_reqId_bits(l2Cache_io_cache_coreResps_3_reqId_bits),
    .io_cache_coreResps_3_rData(l2Cache_io_cache_coreResps_3_rData),
    .io_cache_coreResps_3_responseStatus(l2Cache_io_cache_coreResps_3_responseStatus),
    .io_mem_rChannel_rAddr_ready(l2Cache_io_mem_rChannel_rAddr_ready),
    .io_mem_rChannel_rAddr_valid(l2Cache_io_mem_rChannel_rAddr_valid),
    .io_mem_rChannel_rAddr_bits(l2Cache_io_mem_rChannel_rAddr_bits),
    .io_mem_rChannel_rData_ready(l2Cache_io_mem_rChannel_rData_ready),
    .io_mem_rChannel_rData_valid(l2Cache_io_mem_rChannel_rData_valid),
    .io_mem_rChannel_rData_bits(l2Cache_io_mem_rChannel_rData_bits),
    .io_mem_rChannel_rLast(l2Cache_io_mem_rChannel_rLast),
    .io_mem_wChannel_wAddr_ready(l2Cache_io_mem_wChannel_wAddr_ready),
    .io_mem_wChannel_wAddr_valid(l2Cache_io_mem_wChannel_wAddr_valid),
    .io_mem_wChannel_wAddr_bits(l2Cache_io_mem_wChannel_wAddr_bits),
    .io_mem_wChannel_wData_ready(l2Cache_io_mem_wChannel_wData_ready),
    .io_mem_wChannel_wData_valid(l2Cache_io_mem_wChannel_wData_valid),
    .io_mem_wChannel_wData_bits(l2Cache_io_mem_wChannel_wData_bits),
    .io_mem_wChannel_wLast(l2Cache_io_mem_wChannel_wLast)
  );
  DummyMemory memory ( // @[SharedPipelinedCacheTestTopDe2115.scala 51:22]
    .clock(memory_clock),
    .reset(memory_reset),
    .io_rChannel_rAddr_ready(memory_io_rChannel_rAddr_ready),
    .io_rChannel_rAddr_valid(memory_io_rChannel_rAddr_valid),
    .io_rChannel_rAddr_bits(memory_io_rChannel_rAddr_bits),
    .io_rChannel_rData_ready(memory_io_rChannel_rData_ready),
    .io_rChannel_rData_valid(memory_io_rChannel_rData_valid),
    .io_rChannel_rData_bits(memory_io_rChannel_rData_bits),
    .io_rChannel_rLast(memory_io_rChannel_rLast),
    .io_wChannel_wAddr_ready(memory_io_wChannel_wAddr_ready),
    .io_wChannel_wAddr_valid(memory_io_wChannel_wAddr_valid),
    .io_wChannel_wAddr_bits(memory_io_wChannel_wAddr_bits),
    .io_wChannel_wData_ready(memory_io_wChannel_wData_ready),
    .io_wChannel_wData_valid(memory_io_wChannel_wData_valid),
    .io_wChannel_wData_bits(memory_io_wChannel_wData_bits),
    .io_wChannel_wLast(memory_io_wChannel_wLast)
  );
  assign io_txd = cacheReqCtrl_io_txd; // @[SharedPipelinedCacheTestTopDe2115.scala 87:10]
  assign cacheReqCtrl_clock = clock;
  assign cacheReqCtrl_reset = reset;
  assign cacheReqCtrl_io_rxd = io_rxd; // @[SharedPipelinedCacheTestTopDe2115.scala 86:10]
  assign cacheReqCtrl_io_cache_coreReqs_0_reqId_ready = l2Cache_io_cache_coreReqs_0_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreReqs_1_reqId_ready = l2Cache_io_cache_coreReqs_1_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreReqs_2_reqId_ready = l2Cache_io_cache_coreReqs_2_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreReqs_3_reqId_ready = l2Cache_io_cache_coreReqs_3_reqId_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_0_reqId_valid = l2Cache_io_cache_coreResps_0_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_0_reqId_bits = l2Cache_io_cache_coreResps_0_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_0_rData = l2Cache_io_cache_coreResps_0_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_0_responseStatus = l2Cache_io_cache_coreResps_0_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_1_reqId_valid = l2Cache_io_cache_coreResps_1_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_1_reqId_bits = l2Cache_io_cache_coreResps_1_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_1_rData = l2Cache_io_cache_coreResps_1_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_1_responseStatus = l2Cache_io_cache_coreResps_1_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_2_reqId_valid = l2Cache_io_cache_coreResps_2_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_2_reqId_bits = l2Cache_io_cache_coreResps_2_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_2_rData = l2Cache_io_cache_coreResps_2_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_2_responseStatus = l2Cache_io_cache_coreResps_2_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_3_reqId_valid = l2Cache_io_cache_coreResps_3_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_3_reqId_bits = l2Cache_io_cache_coreResps_3_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_3_rData = l2Cache_io_cache_coreResps_3_rData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign cacheReqCtrl_io_cache_coreResps_3_responseStatus = l2Cache_io_cache_coreResps_3_responseStatus; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_clock = clock;
  assign l2Cache_reset = reset;
  assign l2Cache_io_cache_coreReqs_0_reqId_valid = cacheReqCtrl_io_cache_coreReqs_0_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_0_reqId_bits = cacheReqCtrl_io_cache_coreReqs_0_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_0_addr = cacheReqCtrl_io_cache_coreReqs_0_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_0_rw = cacheReqCtrl_io_cache_coreReqs_0_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_0_wData = cacheReqCtrl_io_cache_coreReqs_0_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_1_reqId_valid = cacheReqCtrl_io_cache_coreReqs_1_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_1_reqId_bits = cacheReqCtrl_io_cache_coreReqs_1_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_1_addr = cacheReqCtrl_io_cache_coreReqs_1_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_1_rw = cacheReqCtrl_io_cache_coreReqs_1_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_1_wData = cacheReqCtrl_io_cache_coreReqs_1_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_2_reqId_valid = cacheReqCtrl_io_cache_coreReqs_2_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_2_reqId_bits = cacheReqCtrl_io_cache_coreReqs_2_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_2_addr = cacheReqCtrl_io_cache_coreReqs_2_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_2_rw = cacheReqCtrl_io_cache_coreReqs_2_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_2_wData = cacheReqCtrl_io_cache_coreReqs_2_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_3_reqId_valid = cacheReqCtrl_io_cache_coreReqs_3_reqId_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_3_reqId_bits = cacheReqCtrl_io_cache_coreReqs_3_reqId_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_3_addr = cacheReqCtrl_io_cache_coreReqs_3_addr; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_3_rw = cacheReqCtrl_io_cache_coreReqs_3_rw; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_cache_coreReqs_3_wData = cacheReqCtrl_io_cache_coreReqs_3_wData; // @[SharedPipelinedCacheTestTopDe2115.scala 60:20]
  assign l2Cache_io_mem_rChannel_rAddr_ready = memory_io_rChannel_rAddr_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 72:39]
  assign l2Cache_io_mem_rChannel_rData_valid = memory_io_rChannel_rData_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 80:28]
  assign l2Cache_io_mem_rChannel_rData_bits = memory_io_rChannel_rData_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 80:28]
  assign l2Cache_io_mem_rChannel_rLast = memory_io_rChannel_rLast; // @[SharedPipelinedCacheTestTopDe2115.scala 81:28]
  assign l2Cache_io_mem_wChannel_wAddr_ready = memory_io_wChannel_wAddr_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 77:39]
  assign l2Cache_io_mem_wChannel_wData_ready = memory_io_wChannel_wData_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 82:28]
  assign memory_clock = clock;
  assign memory_reset = reset;
  assign memory_io_rChannel_rAddr_valid = l2Cache_io_mem_rChannel_rAddr_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 70:34]
  assign memory_io_rChannel_rAddr_bits = l2Cache_io_mem_rChannel_rAddr_bits[14:1]; // @[SharedPipelinedCacheTestTopDe2115.scala 71:70]
  assign memory_io_rChannel_rData_ready = l2Cache_io_mem_rChannel_rData_ready; // @[SharedPipelinedCacheTestTopDe2115.scala 80:28]
  assign memory_io_wChannel_wAddr_valid = l2Cache_io_mem_wChannel_wAddr_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 75:34]
  assign memory_io_wChannel_wAddr_bits = l2Cache_io_mem_wChannel_wAddr_bits[14:1]; // @[SharedPipelinedCacheTestTopDe2115.scala 76:70]
  assign memory_io_wChannel_wData_valid = l2Cache_io_mem_wChannel_wData_valid; // @[SharedPipelinedCacheTestTopDe2115.scala 82:28]
  assign memory_io_wChannel_wData_bits = l2Cache_io_mem_wChannel_wData_bits; // @[SharedPipelinedCacheTestTopDe2115.scala 82:28]
  assign memory_io_wChannel_wLast = l2Cache_io_mem_wChannel_wLast; // @[SharedPipelinedCacheTestTopDe2115.scala 83:28]
endmodule